`timescale 1ns/100ps
module MuxN_2(
    input [54:0] io_ins_9_x,
    input [54:0] io_ins_8_x,
    input [54:0] io_ins_7_x,
    input [54:0] io_ins_6_x,
    input [54:0] io_ins_5_x,
    input [54:0] io_ins_4_x,
    input [54:0] io_ins_3_x,
    input [54:0] io_ins_2_x,
    input [54:0] io_ins_1_x,
    input [54:0] io_ins_0_x,
    input [3:0] io_sel,
    output[54:0] io_out_x
);

  wire[54:0] T0;
  wire[54:0] T1;
  wire[54:0] T2;
  wire[54:0] T3;
  wire T4;
  wire[3:0] T5;
  wire[54:0] T6;
  wire T7;
  wire T8;
  wire[54:0] T9;
  wire[54:0] T10;
  wire T11;
  wire[54:0] T12;
  wire T13;
  wire T14;
  wire T15;
  wire[54:0] T16;
  wire T17;
  wire T18;


  assign io_out_x = T0;
  assign T0 = T18 ? T16 : T1;
  assign T1 = T15 ? T9 : T2;
  assign T2 = T8 ? T6 : T3;
  assign T3 = T4 ? io_ins_1_x : io_ins_0_x;
  assign T4 = T5[1'h0:1'h0];
  assign T5 = io_sel;
  assign T6 = T7 ? io_ins_3_x : io_ins_2_x;
  assign T7 = T5[1'h0:1'h0];
  assign T8 = T5[1'h1:1'h1];
  assign T9 = T14 ? T12 : T10;
  assign T10 = T11 ? io_ins_5_x : io_ins_4_x;
  assign T11 = T5[1'h0:1'h0];
  assign T12 = T13 ? io_ins_7_x : io_ins_6_x;
  assign T13 = T5[1'h0:1'h0];
  assign T14 = T5[1'h1:1'h1];
  assign T15 = T5[2'h2:2'h2];
  assign T16 = T17 ? io_ins_9_x : io_ins_8_x;
  assign T17 = T5[1'h0:1'h0];
  assign T18 = T5[2'h3:2'h3];
endmodule

module Switch(
    input [54:0] io_inPorts_9_x,
    input [54:0] io_inPorts_8_x,
    input [54:0] io_inPorts_7_x,
    input [54:0] io_inPorts_6_x,
    input [54:0] io_inPorts_5_x,
    input [54:0] io_inPorts_4_x,
    input [54:0] io_inPorts_3_x,
    input [54:0] io_inPorts_2_x,
    input [54:0] io_inPorts_1_x,
    input [54:0] io_inPorts_0_x,
    output[54:0] io_outPorts_4_x,
    output[54:0] io_outPorts_3_x,
    output[54:0] io_outPorts_2_x,
    output[54:0] io_outPorts_1_x,
    output[54:0] io_outPorts_0_x,
    input [3:0] io_sel_4,
    input [3:0] io_sel_3,
    input [3:0] io_sel_2,
    input [3:0] io_sel_1,
    input [3:0] io_sel_0
);

  wire[54:0] MuxN_io_out_x;
  wire[54:0] MuxN_1_io_out_x;
  wire[54:0] MuxN_2_io_out_x;
  wire[54:0] MuxN_3_io_out_x;
  wire[54:0] MuxN_4_io_out_x;


  assign io_outPorts_0_x = MuxN_io_out_x;
  assign io_outPorts_1_x = MuxN_1_io_out_x;
  assign io_outPorts_2_x = MuxN_2_io_out_x;
  assign io_outPorts_3_x = MuxN_3_io_out_x;
  assign io_outPorts_4_x = MuxN_4_io_out_x;
  MuxN_2 MuxN(
       .io_ins_9_x( io_inPorts_9_x ),
       .io_ins_8_x( io_inPorts_8_x ),
       .io_ins_7_x( io_inPorts_7_x ),
       .io_ins_6_x( io_inPorts_6_x ),
       .io_ins_5_x( io_inPorts_5_x ),
       .io_ins_4_x( io_inPorts_4_x ),
       .io_ins_3_x( io_inPorts_3_x ),
       .io_ins_2_x( io_inPorts_2_x ),
       .io_ins_1_x( io_inPorts_1_x ),
       .io_ins_0_x( io_inPorts_0_x ),
       .io_sel( io_sel_0 ),
       .io_out_x( MuxN_io_out_x )
  );
  MuxN_2 MuxN_1(
       .io_ins_9_x( io_inPorts_9_x ),
       .io_ins_8_x( io_inPorts_8_x ),
       .io_ins_7_x( io_inPorts_7_x ),
       .io_ins_6_x( io_inPorts_6_x ),
       .io_ins_5_x( io_inPorts_5_x ),
       .io_ins_4_x( io_inPorts_4_x ),
       .io_ins_3_x( io_inPorts_3_x ),
       .io_ins_2_x( io_inPorts_2_x ),
       .io_ins_1_x( io_inPorts_1_x ),
       .io_ins_0_x( io_inPorts_0_x ),
       .io_sel( io_sel_1 ),
       .io_out_x( MuxN_1_io_out_x )
  );
  MuxN_2 MuxN_2(
       .io_ins_9_x( io_inPorts_9_x ),
       .io_ins_8_x( io_inPorts_8_x ),
       .io_ins_7_x( io_inPorts_7_x ),
       .io_ins_6_x( io_inPorts_6_x ),
       .io_ins_5_x( io_inPorts_5_x ),
       .io_ins_4_x( io_inPorts_4_x ),
       .io_ins_3_x( io_inPorts_3_x ),
       .io_ins_2_x( io_inPorts_2_x ),
       .io_ins_1_x( io_inPorts_1_x ),
       .io_ins_0_x( io_inPorts_0_x ),
       .io_sel( io_sel_2 ),
       .io_out_x( MuxN_2_io_out_x )
  );
  MuxN_2 MuxN_3(
       .io_ins_9_x( io_inPorts_9_x ),
       .io_ins_8_x( io_inPorts_8_x ),
       .io_ins_7_x( io_inPorts_7_x ),
       .io_ins_6_x( io_inPorts_6_x ),
       .io_ins_5_x( io_inPorts_5_x ),
       .io_ins_4_x( io_inPorts_4_x ),
       .io_ins_3_x( io_inPorts_3_x ),
       .io_ins_2_x( io_inPorts_2_x ),
       .io_ins_1_x( io_inPorts_1_x ),
       .io_ins_0_x( io_inPorts_0_x ),
       .io_sel( io_sel_3 ),
       .io_out_x( MuxN_3_io_out_x )
  );
  MuxN_2 MuxN_4(
       .io_ins_9_x( io_inPorts_9_x ),
       .io_ins_8_x( io_inPorts_8_x ),
       .io_ins_7_x( io_inPorts_7_x ),
       .io_ins_6_x( io_inPorts_6_x ),
       .io_ins_5_x( io_inPorts_5_x ),
       .io_ins_4_x( io_inPorts_4_x ),
       .io_ins_3_x( io_inPorts_3_x ),
       .io_ins_2_x( io_inPorts_2_x ),
       .io_ins_1_x( io_inPorts_1_x ),
       .io_ins_0_x( io_inPorts_0_x ),
       .io_sel( io_sel_4 ),
       .io_out_x( MuxN_4_io_out_x )
  );
endmodule

module RRArbiterPriority(input clk, input reset,
    input  io_requests_9_releaseLock,
    output io_requests_9_grant,
    input  io_requests_9_request,
    input [2:0] io_requests_9_priorityLevel,
    input  io_requests_8_releaseLock,
    output io_requests_8_grant,
    input  io_requests_8_request,
    input [2:0] io_requests_8_priorityLevel,
    input  io_requests_7_releaseLock,
    output io_requests_7_grant,
    input  io_requests_7_request,
    input [2:0] io_requests_7_priorityLevel,
    input  io_requests_6_releaseLock,
    output io_requests_6_grant,
    input  io_requests_6_request,
    input [2:0] io_requests_6_priorityLevel,
    input  io_requests_5_releaseLock,
    output io_requests_5_grant,
    input  io_requests_5_request,
    input [2:0] io_requests_5_priorityLevel,
    input  io_requests_4_releaseLock,
    output io_requests_4_grant,
    input  io_requests_4_request,
    input [2:0] io_requests_4_priorityLevel,
    input  io_requests_3_releaseLock,
    output io_requests_3_grant,
    input  io_requests_3_request,
    input [2:0] io_requests_3_priorityLevel,
    input  io_requests_2_releaseLock,
    output io_requests_2_grant,
    input  io_requests_2_request,
    input [2:0] io_requests_2_priorityLevel,
    input  io_requests_1_releaseLock,
    output io_requests_1_grant,
    input  io_requests_1_request,
    input [2:0] io_requests_1_priorityLevel,
    input  io_requests_0_releaseLock,
    output io_requests_0_grant,
    input  io_requests_0_request,
    input [2:0] io_requests_0_priorityLevel,
    input  io_resource_ready,
    output io_resource_valid,
    output[3:0] io_chosen
);

  wire[3:0] T645;
  wire[2:0] T646;
  wire[1:0] T647;
  wire T648;
  wire[1:0] T649;
  wire[1:0] T650;
  wire[3:0] T651;
  wire[3:0] T652;
  wire[7:0] T653;
  wire[7:0] T654;
  wire[9:0] winGrant;
  wire[9:0] T1;
  wire[9:0] T2;
  reg [9:0] nextGrant;
  wire[9:0] T655;
  wire[9:0] T3;
  wire[9:0] T4;
  wire T5;
  wire T6;
  wire T7;
  wire lockRelease;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire[3:0] T13;
  wire[3:0] nextGrantUInt;
  wire[3:0] T656;
  wire[2:0] T657;
  wire[1:0] T658;
  wire T659;
  wire[1:0] T660;
  wire[1:0] T661;
  wire[3:0] T662;
  wire[3:0] T663;
  wire[7:0] T664;
  wire[7:0] T665;
  wire[1:0] T666;
  wire[3:0] T667;
  wire[1:0] T668;
  wire T669;
  wire T670;
  wire T671;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire[3:0] T32;
  wire[3:0] T33;
  wire T34;
  wire[9:0] requestsBits;
  wire[4:0] T35;
  wire[2:0] T36;
  wire[1:0] T37;
  wire T38;
  wire T39;
  wire T40;
  wire[1:0] T41;
  wire T42;
  wire T43;
  wire[4:0] T44;
  wire[2:0] T45;
  wire[1:0] T46;
  wire T47;
  wire T48;
  wire T49;
  wire[1:0] T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire[3:0] T56;
  wire[3:0] T57;
  wire T58;
  wire T59;
  wire[9:0] T60;
  wire[9:0] winner;
  wire[9:0] T61;
  wire[9:0] T62;
  wire[9:0] T63;
  wire[9:0] T64;
  wire[4:0] T65;
  wire[2:0] T66;
  wire[1:0] T67;
  wire T68;
  wire T69;
  wire T70;
  reg  PArraySorted_0_0;
  wire T672;
  wire T71;
  wire T72;
  wire T73;
  wire T74;
  wire T75;
  wire T76;
  reg  PArraySorted_1_0;
  wire T673;
  wire T77;
  wire T78;
  wire T79;
  wire T80;
  wire T81;
  wire T82;
  wire T83;
  wire[2:0] T84;
  wire[2:0] T674;
  wire[3:0] pmax;
  wire[3:0] T675;
  wire[2:0] T85;
  wire[2:0] T86;
  wire[2:0] T87;
  wire[2:0] T88;
  wire[2:0] T89;
  wire[2:0] T90;
  wire[2:0] T91;
  wire[2:0] T92;
  wire[2:0] T93;
  wire[2:0] T94;
  wire[2:0] T676;
  wire[1:0] T95;
  wire[1:0] T96;
  wire[1:0] T97;
  wire[1:0] T98;
  wire[1:0] T99;
  wire[1:0] T100;
  wire[1:0] T101;
  wire[1:0] T102;
  wire[1:0] T103;
  wire[1:0] T104;
  wire[1:0] T105;
  wire[1:0] T106;
  wire[1:0] T107;
  wire[1:0] T108;
  wire[1:0] T109;
  wire[1:0] T110;
  wire[1:0] T111;
  wire[1:0] T112;
  wire[1:0] T113;
  wire[1:0] T114;
  wire[1:0] T677;
  wire T115;
  wire T116;
  wire T117;
  wire T118;
  wire T119;
  wire T120;
  wire T121;
  wire T122;
  wire T123;
  wire T124;
  wire T125;
  wire T126;
  wire T127;
  reg  PArraySorted_1_1;
  wire T678;
  wire T128;
  wire T129;
  wire T130;
  wire T131;
  wire T132;
  wire T133;
  wire T134;
  wire T135;
  reg  PArraySorted_1_2;
  wire T679;
  wire T136;
  wire T137;
  wire T138;
  wire T139;
  wire T140;
  wire T141;
  wire T142;
  wire T143;
  reg  PArraySorted_1_3;
  wire T680;
  wire T144;
  wire T145;
  wire T146;
  wire T147;
  wire T148;
  wire T149;
  wire T150;
  wire T151;
  reg  PArraySorted_1_4;
  wire T681;
  wire T152;
  wire T153;
  wire T154;
  wire T155;
  wire T156;
  wire T157;
  wire T158;
  wire T159;
  reg  PArraySorted_1_5;
  wire T682;
  wire T160;
  wire T161;
  wire T162;
  wire T163;
  wire T164;
  wire T165;
  wire T166;
  wire T167;
  reg  PArraySorted_1_6;
  wire T683;
  wire T168;
  wire T169;
  wire T170;
  wire T171;
  wire T172;
  wire T173;
  wire T174;
  wire T175;
  reg  PArraySorted_1_7;
  wire T684;
  wire T176;
  wire T177;
  wire T178;
  wire T179;
  wire T180;
  wire T181;
  wire T182;
  wire T183;
  reg  PArraySorted_1_8;
  wire T685;
  wire T184;
  wire T185;
  wire T186;
  wire T187;
  wire T188;
  wire T189;
  wire T190;
  wire T191;
  reg  PArraySorted_1_9;
  wire T686;
  wire T192;
  wire T193;
  wire T194;
  wire T195;
  wire T196;
  wire T197;
  wire T198;
  wire T199;
  reg  PArraySorted_2_0;
  wire T687;
  wire T200;
  wire T201;
  wire T202;
  wire T203;
  wire T204;
  wire T205;
  wire T206;
  wire T207;
  reg  PArraySorted_2_1;
  wire T688;
  wire T208;
  wire T209;
  wire T210;
  wire T211;
  wire T212;
  wire T213;
  wire T214;
  wire T215;
  reg  PArraySorted_2_2;
  wire T689;
  wire T216;
  wire T217;
  wire T218;
  wire T219;
  wire T220;
  wire T221;
  wire T222;
  wire T223;
  reg  PArraySorted_2_3;
  wire T690;
  wire T224;
  wire T225;
  wire T226;
  wire T227;
  wire T228;
  wire T229;
  wire T230;
  wire T231;
  reg  PArraySorted_2_4;
  wire T691;
  wire T232;
  wire T233;
  wire T234;
  wire T235;
  wire T236;
  wire T237;
  wire T238;
  wire T239;
  reg  PArraySorted_2_5;
  wire T692;
  wire T240;
  wire T241;
  wire T242;
  wire T243;
  wire T244;
  wire T245;
  wire T246;
  wire T247;
  reg  PArraySorted_2_6;
  wire T693;
  wire T248;
  wire T249;
  wire T250;
  wire T251;
  wire T252;
  wire T253;
  wire T254;
  wire T255;
  reg  PArraySorted_2_7;
  wire T694;
  wire T256;
  wire T257;
  wire T258;
  wire T259;
  wire T260;
  wire T261;
  wire T262;
  wire T263;
  reg  PArraySorted_2_8;
  wire T695;
  wire T264;
  wire T265;
  wire T266;
  wire T267;
  wire T268;
  wire T269;
  wire T270;
  wire T271;
  reg  PArraySorted_2_9;
  wire T696;
  wire T272;
  wire T273;
  wire T274;
  wire T275;
  wire T276;
  wire T277;
  wire T278;
  wire T279;
  reg  PArraySorted_3_0;
  wire T697;
  wire T280;
  wire T281;
  wire T282;
  wire T283;
  wire T284;
  wire T285;
  wire T286;
  wire T287;
  reg  PArraySorted_3_1;
  wire T698;
  wire T288;
  wire T289;
  wire T290;
  wire T291;
  wire T292;
  wire T293;
  wire T294;
  wire T295;
  reg  PArraySorted_3_2;
  wire T699;
  wire T296;
  wire T297;
  wire T298;
  wire T299;
  wire T300;
  wire T301;
  wire T302;
  wire T303;
  reg  PArraySorted_3_3;
  wire T700;
  wire T304;
  wire T305;
  wire T306;
  wire T307;
  wire T308;
  wire T309;
  wire T310;
  wire T311;
  reg  PArraySorted_3_4;
  wire T701;
  wire T312;
  wire T313;
  wire T314;
  wire T315;
  wire T316;
  wire T317;
  wire T318;
  wire T319;
  reg  PArraySorted_3_5;
  wire T702;
  wire T320;
  wire T321;
  wire T322;
  wire T323;
  wire T324;
  wire T325;
  wire T326;
  wire T327;
  reg  PArraySorted_3_6;
  wire T703;
  wire T328;
  wire T329;
  wire T330;
  wire T331;
  wire T332;
  wire T333;
  wire T334;
  wire T335;
  reg  PArraySorted_3_7;
  wire T704;
  wire T336;
  wire T337;
  wire T338;
  wire T339;
  wire T340;
  wire T341;
  wire T342;
  wire T343;
  reg  PArraySorted_3_8;
  wire T705;
  wire T344;
  wire T345;
  wire T346;
  wire T347;
  wire T348;
  wire T349;
  wire T350;
  wire T351;
  reg  PArraySorted_3_9;
  wire T706;
  wire T352;
  wire T353;
  wire T354;
  wire T355;
  wire T356;
  wire T357;
  wire T358;
  wire T359;
  wire T360;
  wire T361;
  reg  PArraySorted_4_1;
  wire T707;
  wire T362;
  wire T363;
  wire T364;
  wire T365;
  wire T366;
  wire T367;
  wire T368;
  wire T369;
  reg  PArraySorted_4_2;
  wire T708;
  wire T370;
  wire T371;
  wire T372;
  wire T373;
  wire T374;
  wire T375;
  wire T376;
  wire T377;
  reg  PArraySorted_4_3;
  wire T709;
  wire T378;
  wire T379;
  wire T380;
  wire T381;
  wire T382;
  wire T383;
  wire T384;
  wire T385;
  reg  PArraySorted_4_4;
  wire T710;
  wire T386;
  wire T387;
  wire T388;
  wire T389;
  wire T390;
  wire T391;
  wire T392;
  wire T393;
  reg  PArraySorted_4_5;
  wire T711;
  wire T394;
  wire T395;
  wire T396;
  wire T397;
  wire T398;
  wire T399;
  wire T400;
  wire T401;
  reg  PArraySorted_4_6;
  wire T712;
  wire T402;
  wire T403;
  wire T404;
  wire T405;
  wire T406;
  wire T407;
  wire T408;
  wire T409;
  reg  PArraySorted_4_7;
  wire T713;
  wire T410;
  wire T411;
  wire T412;
  wire T413;
  wire T414;
  wire T415;
  wire T416;
  wire T417;
  reg  PArraySorted_4_8;
  wire T714;
  wire T418;
  wire T419;
  wire T420;
  wire T421;
  wire T422;
  wire T423;
  wire T424;
  wire T425;
  reg  PArraySorted_4_9;
  wire T715;
  wire T426;
  wire T427;
  wire T428;
  wire T429;
  wire T430;
  wire T431;
  wire T432;
  wire T433;
  wire T434;
  reg  PArraySorted_4_0;
  wire T716;
  wire T435;
  wire T436;
  wire T437;
  wire T438;
  wire T439;
  wire T440;
  wire T441;
  wire T442;
  wire T443;
  wire T444;
  reg  PArraySorted_0_1;
  wire T717;
  wire T445;
  wire T446;
  wire T447;
  wire T448;
  wire T449;
  wire T450;
  wire T451;
  wire T452;
  wire T453;
  wire T454;
  wire T455;
  wire T456;
  wire T457;
  wire T458;
  reg  PArraySorted_0_2;
  wire T718;
  wire T459;
  wire T460;
  wire T461;
  wire T462;
  wire T463;
  wire T464;
  wire T465;
  wire T466;
  wire T467;
  wire T468;
  wire T469;
  wire[1:0] T470;
  wire T471;
  wire T472;
  wire T473;
  reg  PArraySorted_0_3;
  wire T719;
  wire T474;
  wire T475;
  wire T476;
  wire T477;
  wire T478;
  wire T479;
  wire T480;
  wire T481;
  wire T482;
  wire T483;
  wire T484;
  wire T485;
  wire T486;
  wire T487;
  reg  PArraySorted_0_4;
  wire T720;
  wire T488;
  wire T489;
  wire T490;
  wire T491;
  wire T492;
  wire T493;
  wire T494;
  wire T495;
  wire T496;
  wire T497;
  wire T498;
  wire[4:0] T499;
  wire[2:0] T500;
  wire[1:0] T501;
  wire T502;
  wire T503;
  wire T504;
  reg  PArraySorted_0_5;
  wire T721;
  wire T505;
  wire T506;
  wire T507;
  wire T508;
  wire T509;
  wire T510;
  wire T511;
  wire T512;
  wire T513;
  wire T514;
  wire T515;
  wire T516;
  wire T517;
  wire T518;
  reg  PArraySorted_0_6;
  wire T722;
  wire T519;
  wire T520;
  wire T521;
  wire T522;
  wire T523;
  wire T524;
  wire T525;
  wire T526;
  wire T527;
  wire T528;
  wire T529;
  wire T530;
  wire T531;
  wire T532;
  reg  PArraySorted_0_7;
  wire T723;
  wire T533;
  wire T534;
  wire T535;
  wire T536;
  wire T537;
  wire T538;
  wire T539;
  wire T540;
  wire T541;
  wire T542;
  wire T543;
  wire[1:0] T544;
  wire T545;
  wire T546;
  wire T547;
  reg  PArraySorted_0_8;
  wire T724;
  wire T548;
  wire T549;
  wire T550;
  wire T551;
  wire T552;
  wire T553;
  wire T554;
  wire T555;
  wire T556;
  wire T557;
  wire T558;
  wire T559;
  wire T560;
  wire T561;
  reg  PArraySorted_0_9;
  wire T725;
  wire T562;
  wire T563;
  wire T564;
  wire T565;
  wire T566;
  wire T567;
  wire T568;
  wire T569;
  wire T570;
  wire T571;
  wire T572;
  wire[9:0] T573;
  wire[9:0] T574;
  wire[10:0] passSelectL0;
  wire[10:0] T575;
  wire[10:0] T576;
  wire[10:0] T577;
  wire[9:0] T578;
  wire T579;
  wire[8:0] T580;
  wire T581;
  wire[10:0] T582;
  wire[9:0] T583;
  wire[9:0] T584;
  wire T585;
  wire[9:0] passSelectL1;
  wire[9:0] T586;
  wire[9:0] T587;
  wire[9:0] T726;
  wire T588;
  wire[9:0] T589;
  wire[9:0] T590;
  wire T591;
  wire T592;
  wire T593;
  wire T594;
  wire[1:0] T727;
  wire[3:0] T728;
  wire[1:0] T729;
  wire T730;
  wire T731;
  wire T732;
  wire T595;
  wire T596;
  wire T597;
  wire T598;
  wire T599;
  wire T600;
  wire[3:0] T601;
  wire T602;
  wire T603;
  wire T604;
  wire T605;
  wire T606;
  wire T607;
  wire T608;
  wire T609;
  wire T610;
  wire T611;
  wire T612;
  wire T613;
  wire T614;
  wire T615;
  wire T616;
  wire T617;
  wire T618;
  wire T619;
  wire T620;
  wire T621;
  wire T622;
  wire T623;
  wire T624;
  wire T625;
  wire T626;
  wire T627;
  wire T628;
  wire T629;
  wire T630;
  wire T631;
  wire T632;
  wire T633;
  wire T634;
  wire T635;
  wire T636;
  wire T637;
  wire T638;
  wire T639;
  wire T640;
  wire T641;
  wire T642;
  wire T643;
  wire T644;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    nextGrant = {1{1'b0}};
    PArraySorted_0_0 = {1{1'b0}};
    PArraySorted_1_0 = {1{1'b0}};
    PArraySorted_1_1 = {1{1'b0}};
    PArraySorted_1_2 = {1{1'b0}};
    PArraySorted_1_3 = {1{1'b0}};
    PArraySorted_1_4 = {1{1'b0}};
    PArraySorted_1_5 = {1{1'b0}};
    PArraySorted_1_6 = {1{1'b0}};
    PArraySorted_1_7 = {1{1'b0}};
    PArraySorted_1_8 = {1{1'b0}};
    PArraySorted_1_9 = {1{1'b0}};
    PArraySorted_2_0 = {1{1'b0}};
    PArraySorted_2_1 = {1{1'b0}};
    PArraySorted_2_2 = {1{1'b0}};
    PArraySorted_2_3 = {1{1'b0}};
    PArraySorted_2_4 = {1{1'b0}};
    PArraySorted_2_5 = {1{1'b0}};
    PArraySorted_2_6 = {1{1'b0}};
    PArraySorted_2_7 = {1{1'b0}};
    PArraySorted_2_8 = {1{1'b0}};
    PArraySorted_2_9 = {1{1'b0}};
    PArraySorted_3_0 = {1{1'b0}};
    PArraySorted_3_1 = {1{1'b0}};
    PArraySorted_3_2 = {1{1'b0}};
    PArraySorted_3_3 = {1{1'b0}};
    PArraySorted_3_4 = {1{1'b0}};
    PArraySorted_3_5 = {1{1'b0}};
    PArraySorted_3_6 = {1{1'b0}};
    PArraySorted_3_7 = {1{1'b0}};
    PArraySorted_3_8 = {1{1'b0}};
    PArraySorted_3_9 = {1{1'b0}};
    PArraySorted_4_1 = {1{1'b0}};
    PArraySorted_4_2 = {1{1'b0}};
    PArraySorted_4_3 = {1{1'b0}};
    PArraySorted_4_4 = {1{1'b0}};
    PArraySorted_4_5 = {1{1'b0}};
    PArraySorted_4_6 = {1{1'b0}};
    PArraySorted_4_7 = {1{1'b0}};
    PArraySorted_4_8 = {1{1'b0}};
    PArraySorted_4_9 = {1{1'b0}};
    PArraySorted_4_0 = {1{1'b0}};
    PArraySorted_0_1 = {1{1'b0}};
    PArraySorted_0_2 = {1{1'b0}};
    PArraySorted_0_3 = {1{1'b0}};
    PArraySorted_0_4 = {1{1'b0}};
    PArraySorted_0_5 = {1{1'b0}};
    PArraySorted_0_6 = {1{1'b0}};
    PArraySorted_0_7 = {1{1'b0}};
    PArraySorted_0_8 = {1{1'b0}};
    PArraySorted_0_9 = {1{1'b0}};
  end
// synthesis translate_on
`endif

  assign io_chosen = T645;
  assign T645 = {T732, T646};
  assign T646 = {T731, T647};
  assign T647 = {T730, T648};
  assign T648 = T649[1'h1:1'h1];
  assign T649 = T729 | T650;
  assign T650 = T651[1'h1:1'h0];
  assign T651 = T728 | T652;
  assign T652 = T653[2'h3:1'h0];
  assign T653 = T727 | T654;
  assign T654 = winGrant[3'h7:1'h0];
  assign winGrant = T1;
  assign T1 = T593 ? T60 : T2;
  assign T2 = T5 ? nextGrant : 10'h200;
  assign T655 = reset ? 10'h200 : T3;
  assign T3 = T593 ? winGrant : T4;
  assign T4 = T5 ? winGrant : nextGrant;
  assign T5 = T59 & T6;
  assign T6 = T28 & T7;
  assign T7 = ~ lockRelease;
  assign lockRelease = T8;
  assign T8 = T27 ? T25 : T9;
  assign T9 = T24 ? T18 : T10;
  assign T10 = T17 ? T15 : T11;
  assign T11 = T12 ? io_requests_1_releaseLock : io_requests_0_releaseLock;
  assign T12 = T13[1'h0:1'h0];
  assign T13 = nextGrantUInt;
  assign nextGrantUInt = T656;
  assign T656 = {T671, T657};
  assign T657 = {T670, T658};
  assign T658 = {T669, T659};
  assign T659 = T660[1'h1:1'h1];
  assign T660 = T668 | T661;
  assign T661 = T662[1'h1:1'h0];
  assign T662 = T667 | T663;
  assign T663 = T664[2'h3:1'h0];
  assign T664 = T666 | T665;
  assign T665 = nextGrant[3'h7:1'h0];
  assign T666 = nextGrant[4'h9:4'h8];
  assign T667 = T664[3'h7:3'h4];
  assign T668 = T662[2'h3:2'h2];
  assign T669 = T668 != 2'h0;
  assign T670 = T667 != 4'h0;
  assign T671 = T666 != 2'h0;
  assign T15 = T16 ? io_requests_3_releaseLock : io_requests_2_releaseLock;
  assign T16 = T13[1'h0:1'h0];
  assign T17 = T13[1'h1:1'h1];
  assign T18 = T23 ? T21 : T19;
  assign T19 = T20 ? io_requests_5_releaseLock : io_requests_4_releaseLock;
  assign T20 = T13[1'h0:1'h0];
  assign T21 = T22 ? io_requests_7_releaseLock : io_requests_6_releaseLock;
  assign T22 = T13[1'h0:1'h0];
  assign T23 = T13[1'h1:1'h1];
  assign T24 = T13[2'h2:2'h2];
  assign T25 = T26 ? io_requests_9_releaseLock : io_requests_8_releaseLock;
  assign T26 = T13[1'h0:1'h0];
  assign T27 = T13[2'h3:2'h3];
  assign T28 = T53 & T29;
  assign T29 = T34 & T30;
  assign T30 = T31 - 1'h1;
  assign T31 = 1'h1 << T32;
  assign T32 = T33 + 4'h1;
  assign T33 = nextGrantUInt - nextGrantUInt;
  assign T34 = requestsBits >> nextGrantUInt;
  assign requestsBits = {T44, T35};
  assign T35 = {T41, T36};
  assign T36 = {T40, T37};
  assign T37 = {T39, T38};
  assign T38 = io_requests_0_request;
  assign T39 = io_requests_1_request;
  assign T40 = io_requests_2_request;
  assign T41 = {T43, T42};
  assign T42 = io_requests_3_request;
  assign T43 = io_requests_4_request;
  assign T44 = {T50, T45};
  assign T45 = {T49, T46};
  assign T46 = {T48, T47};
  assign T47 = io_requests_5_request;
  assign T48 = io_requests_6_request;
  assign T49 = io_requests_7_request;
  assign T50 = {T52, T51};
  assign T51 = io_requests_8_request;
  assign T52 = io_requests_9_request;
  assign T53 = T58 & T54;
  assign T54 = T55 - 1'h1;
  assign T55 = 1'h1 << T56;
  assign T56 = T57 + 4'h1;
  assign T57 = nextGrantUInt - nextGrantUInt;
  assign T58 = nextGrant >> nextGrantUInt;
  assign T59 = requestsBits != 10'h0;
  assign T60 = T592 ? winner : nextGrant;
  assign winner = T61;
  assign T61 = T593 ? T62 : 10'h0;
  assign T62 = T573 & T63;
  assign T63 = T64;
  assign T64 = {T499, T65};
  assign T65 = {T470, T66};
  assign T66 = {T456, T67};
  assign T67 = {T442, T68};
  assign T68 = T441 ? PArraySorted_4_0 : T69;
  assign T69 = T434 ? T432 : T70;
  assign T70 = T83 ? PArraySorted_1_0 : PArraySorted_0_0;
  assign T672 = reset ? 1'h0 : T71;
  assign T71 = T73 ? 1'h1 : T72;
  assign T72 = T593 ? 1'h0 : PArraySorted_0_0;
  assign T73 = T75 & T74;
  assign T74 = requestsBits[1'h0:1'h0];
  assign T75 = T593 & T76;
  assign T76 = io_requests_0_priorityLevel == 3'h0;
  assign T673 = reset ? 1'h0 : T77;
  assign T77 = T79 ? 1'h1 : T78;
  assign T78 = T593 ? 1'h0 : PArraySorted_1_0;
  assign T79 = T81 & T80;
  assign T80 = requestsBits[1'h0:1'h0];
  assign T81 = T593 & T82;
  assign T82 = io_requests_0_priorityLevel == 3'h1;
  assign T83 = T84[1'h0:1'h0];
  assign T84 = T674;
  assign T674 = pmax[2'h2:1'h0];
  assign pmax = T675;
  assign T675 = {1'h0, T85};
  assign T85 = T424 ? 3'h4 : T86;
  assign T86 = T416 ? 3'h4 : T87;
  assign T87 = T408 ? 3'h4 : T88;
  assign T88 = T400 ? 3'h4 : T89;
  assign T89 = T392 ? 3'h4 : T90;
  assign T90 = T384 ? 3'h4 : T91;
  assign T91 = T376 ? 3'h4 : T92;
  assign T92 = T368 ? 3'h4 : T93;
  assign T93 = T360 ? 3'h4 : T94;
  assign T94 = T358 ? 3'h4 : T676;
  assign T676 = {1'h0, T95};
  assign T95 = T350 ? 2'h3 : T96;
  assign T96 = T342 ? 2'h3 : T97;
  assign T97 = T334 ? 2'h3 : T98;
  assign T98 = T326 ? 2'h3 : T99;
  assign T99 = T318 ? 2'h3 : T100;
  assign T100 = T310 ? 2'h3 : T101;
  assign T101 = T302 ? 2'h3 : T102;
  assign T102 = T294 ? 2'h3 : T103;
  assign T103 = T286 ? 2'h3 : T104;
  assign T104 = T278 ? 2'h3 : T105;
  assign T105 = T270 ? 2'h2 : T106;
  assign T106 = T262 ? 2'h2 : T107;
  assign T107 = T254 ? 2'h2 : T108;
  assign T108 = T246 ? 2'h2 : T109;
  assign T109 = T238 ? 2'h2 : T110;
  assign T110 = T230 ? 2'h2 : T111;
  assign T111 = T222 ? 2'h2 : T112;
  assign T112 = T214 ? 2'h2 : T113;
  assign T113 = T206 ? 2'h2 : T114;
  assign T114 = T198 ? 2'h2 : T677;
  assign T677 = {1'h0, T115};
  assign T115 = T190 ? 1'h1 : T116;
  assign T116 = T182 ? 1'h1 : T117;
  assign T117 = T174 ? 1'h1 : T118;
  assign T118 = T166 ? 1'h1 : T119;
  assign T119 = T158 ? 1'h1 : T120;
  assign T120 = T150 ? 1'h1 : T121;
  assign T121 = T142 ? 1'h1 : T122;
  assign T122 = T134 ? 1'h1 : T123;
  assign T123 = T126 ? 1'h1 : T124;
  assign T124 = T593 & T125;
  assign T125 = PArraySorted_1_0 == 1'h1;
  assign T126 = T593 & T127;
  assign T127 = PArraySorted_1_1 == 1'h1;
  assign T678 = reset ? 1'h0 : T128;
  assign T128 = T130 ? 1'h1 : T129;
  assign T129 = T593 ? 1'h0 : PArraySorted_1_1;
  assign T130 = T132 & T131;
  assign T131 = requestsBits[1'h1:1'h1];
  assign T132 = T593 & T133;
  assign T133 = io_requests_1_priorityLevel == 3'h1;
  assign T134 = T593 & T135;
  assign T135 = PArraySorted_1_2 == 1'h1;
  assign T679 = reset ? 1'h0 : T136;
  assign T136 = T138 ? 1'h1 : T137;
  assign T137 = T593 ? 1'h0 : PArraySorted_1_2;
  assign T138 = T140 & T139;
  assign T139 = requestsBits[2'h2:2'h2];
  assign T140 = T593 & T141;
  assign T141 = io_requests_2_priorityLevel == 3'h1;
  assign T142 = T593 & T143;
  assign T143 = PArraySorted_1_3 == 1'h1;
  assign T680 = reset ? 1'h0 : T144;
  assign T144 = T146 ? 1'h1 : T145;
  assign T145 = T593 ? 1'h0 : PArraySorted_1_3;
  assign T146 = T148 & T147;
  assign T147 = requestsBits[2'h3:2'h3];
  assign T148 = T593 & T149;
  assign T149 = io_requests_3_priorityLevel == 3'h1;
  assign T150 = T593 & T151;
  assign T151 = PArraySorted_1_4 == 1'h1;
  assign T681 = reset ? 1'h0 : T152;
  assign T152 = T154 ? 1'h1 : T153;
  assign T153 = T593 ? 1'h0 : PArraySorted_1_4;
  assign T154 = T156 & T155;
  assign T155 = requestsBits[3'h4:3'h4];
  assign T156 = T593 & T157;
  assign T157 = io_requests_4_priorityLevel == 3'h1;
  assign T158 = T593 & T159;
  assign T159 = PArraySorted_1_5 == 1'h1;
  assign T682 = reset ? 1'h0 : T160;
  assign T160 = T162 ? 1'h1 : T161;
  assign T161 = T593 ? 1'h0 : PArraySorted_1_5;
  assign T162 = T164 & T163;
  assign T163 = requestsBits[3'h5:3'h5];
  assign T164 = T593 & T165;
  assign T165 = io_requests_5_priorityLevel == 3'h1;
  assign T166 = T593 & T167;
  assign T167 = PArraySorted_1_6 == 1'h1;
  assign T683 = reset ? 1'h0 : T168;
  assign T168 = T170 ? 1'h1 : T169;
  assign T169 = T593 ? 1'h0 : PArraySorted_1_6;
  assign T170 = T172 & T171;
  assign T171 = requestsBits[3'h6:3'h6];
  assign T172 = T593 & T173;
  assign T173 = io_requests_6_priorityLevel == 3'h1;
  assign T174 = T593 & T175;
  assign T175 = PArraySorted_1_7 == 1'h1;
  assign T684 = reset ? 1'h0 : T176;
  assign T176 = T178 ? 1'h1 : T177;
  assign T177 = T593 ? 1'h0 : PArraySorted_1_7;
  assign T178 = T180 & T179;
  assign T179 = requestsBits[3'h7:3'h7];
  assign T180 = T593 & T181;
  assign T181 = io_requests_7_priorityLevel == 3'h1;
  assign T182 = T593 & T183;
  assign T183 = PArraySorted_1_8 == 1'h1;
  assign T685 = reset ? 1'h0 : T184;
  assign T184 = T186 ? 1'h1 : T185;
  assign T185 = T593 ? 1'h0 : PArraySorted_1_8;
  assign T186 = T188 & T187;
  assign T187 = requestsBits[4'h8:4'h8];
  assign T188 = T593 & T189;
  assign T189 = io_requests_8_priorityLevel == 3'h1;
  assign T190 = T593 & T191;
  assign T191 = PArraySorted_1_9 == 1'h1;
  assign T686 = reset ? 1'h0 : T192;
  assign T192 = T194 ? 1'h1 : T193;
  assign T193 = T593 ? 1'h0 : PArraySorted_1_9;
  assign T194 = T196 & T195;
  assign T195 = requestsBits[4'h9:4'h9];
  assign T196 = T593 & T197;
  assign T197 = io_requests_9_priorityLevel == 3'h1;
  assign T198 = T593 & T199;
  assign T199 = PArraySorted_2_0 == 1'h1;
  assign T687 = reset ? 1'h0 : T200;
  assign T200 = T202 ? 1'h1 : T201;
  assign T201 = T593 ? 1'h0 : PArraySorted_2_0;
  assign T202 = T204 & T203;
  assign T203 = requestsBits[1'h0:1'h0];
  assign T204 = T593 & T205;
  assign T205 = io_requests_0_priorityLevel == 3'h2;
  assign T206 = T593 & T207;
  assign T207 = PArraySorted_2_1 == 1'h1;
  assign T688 = reset ? 1'h0 : T208;
  assign T208 = T210 ? 1'h1 : T209;
  assign T209 = T593 ? 1'h0 : PArraySorted_2_1;
  assign T210 = T212 & T211;
  assign T211 = requestsBits[1'h1:1'h1];
  assign T212 = T593 & T213;
  assign T213 = io_requests_1_priorityLevel == 3'h2;
  assign T214 = T593 & T215;
  assign T215 = PArraySorted_2_2 == 1'h1;
  assign T689 = reset ? 1'h0 : T216;
  assign T216 = T218 ? 1'h1 : T217;
  assign T217 = T593 ? 1'h0 : PArraySorted_2_2;
  assign T218 = T220 & T219;
  assign T219 = requestsBits[2'h2:2'h2];
  assign T220 = T593 & T221;
  assign T221 = io_requests_2_priorityLevel == 3'h2;
  assign T222 = T593 & T223;
  assign T223 = PArraySorted_2_3 == 1'h1;
  assign T690 = reset ? 1'h0 : T224;
  assign T224 = T226 ? 1'h1 : T225;
  assign T225 = T593 ? 1'h0 : PArraySorted_2_3;
  assign T226 = T228 & T227;
  assign T227 = requestsBits[2'h3:2'h3];
  assign T228 = T593 & T229;
  assign T229 = io_requests_3_priorityLevel == 3'h2;
  assign T230 = T593 & T231;
  assign T231 = PArraySorted_2_4 == 1'h1;
  assign T691 = reset ? 1'h0 : T232;
  assign T232 = T234 ? 1'h1 : T233;
  assign T233 = T593 ? 1'h0 : PArraySorted_2_4;
  assign T234 = T236 & T235;
  assign T235 = requestsBits[3'h4:3'h4];
  assign T236 = T593 & T237;
  assign T237 = io_requests_4_priorityLevel == 3'h2;
  assign T238 = T593 & T239;
  assign T239 = PArraySorted_2_5 == 1'h1;
  assign T692 = reset ? 1'h0 : T240;
  assign T240 = T242 ? 1'h1 : T241;
  assign T241 = T593 ? 1'h0 : PArraySorted_2_5;
  assign T242 = T244 & T243;
  assign T243 = requestsBits[3'h5:3'h5];
  assign T244 = T593 & T245;
  assign T245 = io_requests_5_priorityLevel == 3'h2;
  assign T246 = T593 & T247;
  assign T247 = PArraySorted_2_6 == 1'h1;
  assign T693 = reset ? 1'h0 : T248;
  assign T248 = T250 ? 1'h1 : T249;
  assign T249 = T593 ? 1'h0 : PArraySorted_2_6;
  assign T250 = T252 & T251;
  assign T251 = requestsBits[3'h6:3'h6];
  assign T252 = T593 & T253;
  assign T253 = io_requests_6_priorityLevel == 3'h2;
  assign T254 = T593 & T255;
  assign T255 = PArraySorted_2_7 == 1'h1;
  assign T694 = reset ? 1'h0 : T256;
  assign T256 = T258 ? 1'h1 : T257;
  assign T257 = T593 ? 1'h0 : PArraySorted_2_7;
  assign T258 = T260 & T259;
  assign T259 = requestsBits[3'h7:3'h7];
  assign T260 = T593 & T261;
  assign T261 = io_requests_7_priorityLevel == 3'h2;
  assign T262 = T593 & T263;
  assign T263 = PArraySorted_2_8 == 1'h1;
  assign T695 = reset ? 1'h0 : T264;
  assign T264 = T266 ? 1'h1 : T265;
  assign T265 = T593 ? 1'h0 : PArraySorted_2_8;
  assign T266 = T268 & T267;
  assign T267 = requestsBits[4'h8:4'h8];
  assign T268 = T593 & T269;
  assign T269 = io_requests_8_priorityLevel == 3'h2;
  assign T270 = T593 & T271;
  assign T271 = PArraySorted_2_9 == 1'h1;
  assign T696 = reset ? 1'h0 : T272;
  assign T272 = T274 ? 1'h1 : T273;
  assign T273 = T593 ? 1'h0 : PArraySorted_2_9;
  assign T274 = T276 & T275;
  assign T275 = requestsBits[4'h9:4'h9];
  assign T276 = T593 & T277;
  assign T277 = io_requests_9_priorityLevel == 3'h2;
  assign T278 = T593 & T279;
  assign T279 = PArraySorted_3_0 == 1'h1;
  assign T697 = reset ? 1'h0 : T280;
  assign T280 = T282 ? 1'h1 : T281;
  assign T281 = T593 ? 1'h0 : PArraySorted_3_0;
  assign T282 = T284 & T283;
  assign T283 = requestsBits[1'h0:1'h0];
  assign T284 = T593 & T285;
  assign T285 = io_requests_0_priorityLevel == 3'h3;
  assign T286 = T593 & T287;
  assign T287 = PArraySorted_3_1 == 1'h1;
  assign T698 = reset ? 1'h0 : T288;
  assign T288 = T290 ? 1'h1 : T289;
  assign T289 = T593 ? 1'h0 : PArraySorted_3_1;
  assign T290 = T292 & T291;
  assign T291 = requestsBits[1'h1:1'h1];
  assign T292 = T593 & T293;
  assign T293 = io_requests_1_priorityLevel == 3'h3;
  assign T294 = T593 & T295;
  assign T295 = PArraySorted_3_2 == 1'h1;
  assign T699 = reset ? 1'h0 : T296;
  assign T296 = T298 ? 1'h1 : T297;
  assign T297 = T593 ? 1'h0 : PArraySorted_3_2;
  assign T298 = T300 & T299;
  assign T299 = requestsBits[2'h2:2'h2];
  assign T300 = T593 & T301;
  assign T301 = io_requests_2_priorityLevel == 3'h3;
  assign T302 = T593 & T303;
  assign T303 = PArraySorted_3_3 == 1'h1;
  assign T700 = reset ? 1'h0 : T304;
  assign T304 = T306 ? 1'h1 : T305;
  assign T305 = T593 ? 1'h0 : PArraySorted_3_3;
  assign T306 = T308 & T307;
  assign T307 = requestsBits[2'h3:2'h3];
  assign T308 = T593 & T309;
  assign T309 = io_requests_3_priorityLevel == 3'h3;
  assign T310 = T593 & T311;
  assign T311 = PArraySorted_3_4 == 1'h1;
  assign T701 = reset ? 1'h0 : T312;
  assign T312 = T314 ? 1'h1 : T313;
  assign T313 = T593 ? 1'h0 : PArraySorted_3_4;
  assign T314 = T316 & T315;
  assign T315 = requestsBits[3'h4:3'h4];
  assign T316 = T593 & T317;
  assign T317 = io_requests_4_priorityLevel == 3'h3;
  assign T318 = T593 & T319;
  assign T319 = PArraySorted_3_5 == 1'h1;
  assign T702 = reset ? 1'h0 : T320;
  assign T320 = T322 ? 1'h1 : T321;
  assign T321 = T593 ? 1'h0 : PArraySorted_3_5;
  assign T322 = T324 & T323;
  assign T323 = requestsBits[3'h5:3'h5];
  assign T324 = T593 & T325;
  assign T325 = io_requests_5_priorityLevel == 3'h3;
  assign T326 = T593 & T327;
  assign T327 = PArraySorted_3_6 == 1'h1;
  assign T703 = reset ? 1'h0 : T328;
  assign T328 = T330 ? 1'h1 : T329;
  assign T329 = T593 ? 1'h0 : PArraySorted_3_6;
  assign T330 = T332 & T331;
  assign T331 = requestsBits[3'h6:3'h6];
  assign T332 = T593 & T333;
  assign T333 = io_requests_6_priorityLevel == 3'h3;
  assign T334 = T593 & T335;
  assign T335 = PArraySorted_3_7 == 1'h1;
  assign T704 = reset ? 1'h0 : T336;
  assign T336 = T338 ? 1'h1 : T337;
  assign T337 = T593 ? 1'h0 : PArraySorted_3_7;
  assign T338 = T340 & T339;
  assign T339 = requestsBits[3'h7:3'h7];
  assign T340 = T593 & T341;
  assign T341 = io_requests_7_priorityLevel == 3'h3;
  assign T342 = T593 & T343;
  assign T343 = PArraySorted_3_8 == 1'h1;
  assign T705 = reset ? 1'h0 : T344;
  assign T344 = T346 ? 1'h1 : T345;
  assign T345 = T593 ? 1'h0 : PArraySorted_3_8;
  assign T346 = T348 & T347;
  assign T347 = requestsBits[4'h8:4'h8];
  assign T348 = T593 & T349;
  assign T349 = io_requests_8_priorityLevel == 3'h3;
  assign T350 = T593 & T351;
  assign T351 = PArraySorted_3_9 == 1'h1;
  assign T706 = reset ? 1'h0 : T352;
  assign T352 = T354 ? 1'h1 : T353;
  assign T353 = T593 ? 1'h0 : PArraySorted_3_9;
  assign T354 = T356 & T355;
  assign T355 = requestsBits[4'h9:4'h9];
  assign T356 = T593 & T357;
  assign T357 = io_requests_9_priorityLevel == 3'h3;
  assign T358 = T593 & T359;
  assign T359 = PArraySorted_4_0 == 1'h1;
  assign T360 = T593 & T361;
  assign T361 = PArraySorted_4_1 == 1'h1;
  assign T707 = reset ? 1'h0 : T362;
  assign T362 = T364 ? 1'h1 : T363;
  assign T363 = T593 ? 1'h0 : PArraySorted_4_1;
  assign T364 = T366 & T365;
  assign T365 = requestsBits[1'h1:1'h1];
  assign T366 = T593 & T367;
  assign T367 = io_requests_1_priorityLevel == 3'h4;
  assign T368 = T593 & T369;
  assign T369 = PArraySorted_4_2 == 1'h1;
  assign T708 = reset ? 1'h0 : T370;
  assign T370 = T372 ? 1'h1 : T371;
  assign T371 = T593 ? 1'h0 : PArraySorted_4_2;
  assign T372 = T374 & T373;
  assign T373 = requestsBits[2'h2:2'h2];
  assign T374 = T593 & T375;
  assign T375 = io_requests_2_priorityLevel == 3'h4;
  assign T376 = T593 & T377;
  assign T377 = PArraySorted_4_3 == 1'h1;
  assign T709 = reset ? 1'h0 : T378;
  assign T378 = T380 ? 1'h1 : T379;
  assign T379 = T593 ? 1'h0 : PArraySorted_4_3;
  assign T380 = T382 & T381;
  assign T381 = requestsBits[2'h3:2'h3];
  assign T382 = T593 & T383;
  assign T383 = io_requests_3_priorityLevel == 3'h4;
  assign T384 = T593 & T385;
  assign T385 = PArraySorted_4_4 == 1'h1;
  assign T710 = reset ? 1'h0 : T386;
  assign T386 = T388 ? 1'h1 : T387;
  assign T387 = T593 ? 1'h0 : PArraySorted_4_4;
  assign T388 = T390 & T389;
  assign T389 = requestsBits[3'h4:3'h4];
  assign T390 = T593 & T391;
  assign T391 = io_requests_4_priorityLevel == 3'h4;
  assign T392 = T593 & T393;
  assign T393 = PArraySorted_4_5 == 1'h1;
  assign T711 = reset ? 1'h0 : T394;
  assign T394 = T396 ? 1'h1 : T395;
  assign T395 = T593 ? 1'h0 : PArraySorted_4_5;
  assign T396 = T398 & T397;
  assign T397 = requestsBits[3'h5:3'h5];
  assign T398 = T593 & T399;
  assign T399 = io_requests_5_priorityLevel == 3'h4;
  assign T400 = T593 & T401;
  assign T401 = PArraySorted_4_6 == 1'h1;
  assign T712 = reset ? 1'h0 : T402;
  assign T402 = T404 ? 1'h1 : T403;
  assign T403 = T593 ? 1'h0 : PArraySorted_4_6;
  assign T404 = T406 & T405;
  assign T405 = requestsBits[3'h6:3'h6];
  assign T406 = T593 & T407;
  assign T407 = io_requests_6_priorityLevel == 3'h4;
  assign T408 = T593 & T409;
  assign T409 = PArraySorted_4_7 == 1'h1;
  assign T713 = reset ? 1'h0 : T410;
  assign T410 = T412 ? 1'h1 : T411;
  assign T411 = T593 ? 1'h0 : PArraySorted_4_7;
  assign T412 = T414 & T413;
  assign T413 = requestsBits[3'h7:3'h7];
  assign T414 = T593 & T415;
  assign T415 = io_requests_7_priorityLevel == 3'h4;
  assign T416 = T593 & T417;
  assign T417 = PArraySorted_4_8 == 1'h1;
  assign T714 = reset ? 1'h0 : T418;
  assign T418 = T420 ? 1'h1 : T419;
  assign T419 = T593 ? 1'h0 : PArraySorted_4_8;
  assign T420 = T422 & T421;
  assign T421 = requestsBits[4'h8:4'h8];
  assign T422 = T593 & T423;
  assign T423 = io_requests_8_priorityLevel == 3'h4;
  assign T424 = T593 & T425;
  assign T425 = PArraySorted_4_9 == 1'h1;
  assign T715 = reset ? 1'h0 : T426;
  assign T426 = T428 ? 1'h1 : T427;
  assign T427 = T593 ? 1'h0 : PArraySorted_4_9;
  assign T428 = T430 & T429;
  assign T429 = requestsBits[4'h9:4'h9];
  assign T430 = T593 & T431;
  assign T431 = io_requests_9_priorityLevel == 3'h4;
  assign T432 = T433 ? PArraySorted_3_0 : PArraySorted_2_0;
  assign T433 = T84[1'h0:1'h0];
  assign T434 = T84[1'h1:1'h1];
  assign T716 = reset ? 1'h0 : T435;
  assign T435 = T437 ? 1'h1 : T436;
  assign T436 = T593 ? 1'h0 : PArraySorted_4_0;
  assign T437 = T439 & T438;
  assign T438 = requestsBits[1'h0:1'h0];
  assign T439 = T593 & T440;
  assign T440 = io_requests_0_priorityLevel == 3'h4;
  assign T441 = T84[2'h2:2'h2];
  assign T442 = T455 ? PArraySorted_4_1 : T443;
  assign T443 = T454 ? T452 : T444;
  assign T444 = T451 ? PArraySorted_1_1 : PArraySorted_0_1;
  assign T717 = reset ? 1'h0 : T445;
  assign T445 = T447 ? 1'h1 : T446;
  assign T446 = T593 ? 1'h0 : PArraySorted_0_1;
  assign T447 = T449 & T448;
  assign T448 = requestsBits[1'h1:1'h1];
  assign T449 = T593 & T450;
  assign T450 = io_requests_1_priorityLevel == 3'h0;
  assign T451 = T84[1'h0:1'h0];
  assign T452 = T453 ? PArraySorted_3_1 : PArraySorted_2_1;
  assign T453 = T84[1'h0:1'h0];
  assign T454 = T84[1'h1:1'h1];
  assign T455 = T84[2'h2:2'h2];
  assign T456 = T469 ? PArraySorted_4_2 : T457;
  assign T457 = T468 ? T466 : T458;
  assign T458 = T465 ? PArraySorted_1_2 : PArraySorted_0_2;
  assign T718 = reset ? 1'h0 : T459;
  assign T459 = T461 ? 1'h1 : T460;
  assign T460 = T593 ? 1'h0 : PArraySorted_0_2;
  assign T461 = T463 & T462;
  assign T462 = requestsBits[2'h2:2'h2];
  assign T463 = T593 & T464;
  assign T464 = io_requests_2_priorityLevel == 3'h0;
  assign T465 = T84[1'h0:1'h0];
  assign T466 = T467 ? PArraySorted_3_2 : PArraySorted_2_2;
  assign T467 = T84[1'h0:1'h0];
  assign T468 = T84[1'h1:1'h1];
  assign T469 = T84[2'h2:2'h2];
  assign T470 = {T485, T471};
  assign T471 = T484 ? PArraySorted_4_3 : T472;
  assign T472 = T483 ? T481 : T473;
  assign T473 = T480 ? PArraySorted_1_3 : PArraySorted_0_3;
  assign T719 = reset ? 1'h0 : T474;
  assign T474 = T476 ? 1'h1 : T475;
  assign T475 = T593 ? 1'h0 : PArraySorted_0_3;
  assign T476 = T478 & T477;
  assign T477 = requestsBits[2'h3:2'h3];
  assign T478 = T593 & T479;
  assign T479 = io_requests_3_priorityLevel == 3'h0;
  assign T480 = T84[1'h0:1'h0];
  assign T481 = T482 ? PArraySorted_3_3 : PArraySorted_2_3;
  assign T482 = T84[1'h0:1'h0];
  assign T483 = T84[1'h1:1'h1];
  assign T484 = T84[2'h2:2'h2];
  assign T485 = T498 ? PArraySorted_4_4 : T486;
  assign T486 = T497 ? T495 : T487;
  assign T487 = T494 ? PArraySorted_1_4 : PArraySorted_0_4;
  assign T720 = reset ? 1'h0 : T488;
  assign T488 = T490 ? 1'h1 : T489;
  assign T489 = T593 ? 1'h0 : PArraySorted_0_4;
  assign T490 = T492 & T491;
  assign T491 = requestsBits[3'h4:3'h4];
  assign T492 = T593 & T493;
  assign T493 = io_requests_4_priorityLevel == 3'h0;
  assign T494 = T84[1'h0:1'h0];
  assign T495 = T496 ? PArraySorted_3_4 : PArraySorted_2_4;
  assign T496 = T84[1'h0:1'h0];
  assign T497 = T84[1'h1:1'h1];
  assign T498 = T84[2'h2:2'h2];
  assign T499 = {T544, T500};
  assign T500 = {T530, T501};
  assign T501 = {T516, T502};
  assign T502 = T515 ? PArraySorted_4_5 : T503;
  assign T503 = T514 ? T512 : T504;
  assign T504 = T511 ? PArraySorted_1_5 : PArraySorted_0_5;
  assign T721 = reset ? 1'h0 : T505;
  assign T505 = T507 ? 1'h1 : T506;
  assign T506 = T593 ? 1'h0 : PArraySorted_0_5;
  assign T507 = T509 & T508;
  assign T508 = requestsBits[3'h5:3'h5];
  assign T509 = T593 & T510;
  assign T510 = io_requests_5_priorityLevel == 3'h0;
  assign T511 = T84[1'h0:1'h0];
  assign T512 = T513 ? PArraySorted_3_5 : PArraySorted_2_5;
  assign T513 = T84[1'h0:1'h0];
  assign T514 = T84[1'h1:1'h1];
  assign T515 = T84[2'h2:2'h2];
  assign T516 = T529 ? PArraySorted_4_6 : T517;
  assign T517 = T528 ? T526 : T518;
  assign T518 = T525 ? PArraySorted_1_6 : PArraySorted_0_6;
  assign T722 = reset ? 1'h0 : T519;
  assign T519 = T521 ? 1'h1 : T520;
  assign T520 = T593 ? 1'h0 : PArraySorted_0_6;
  assign T521 = T523 & T522;
  assign T522 = requestsBits[3'h6:3'h6];
  assign T523 = T593 & T524;
  assign T524 = io_requests_6_priorityLevel == 3'h0;
  assign T525 = T84[1'h0:1'h0];
  assign T526 = T527 ? PArraySorted_3_6 : PArraySorted_2_6;
  assign T527 = T84[1'h0:1'h0];
  assign T528 = T84[1'h1:1'h1];
  assign T529 = T84[2'h2:2'h2];
  assign T530 = T543 ? PArraySorted_4_7 : T531;
  assign T531 = T542 ? T540 : T532;
  assign T532 = T539 ? PArraySorted_1_7 : PArraySorted_0_7;
  assign T723 = reset ? 1'h0 : T533;
  assign T533 = T535 ? 1'h1 : T534;
  assign T534 = T593 ? 1'h0 : PArraySorted_0_7;
  assign T535 = T537 & T536;
  assign T536 = requestsBits[3'h7:3'h7];
  assign T537 = T593 & T538;
  assign T538 = io_requests_7_priorityLevel == 3'h0;
  assign T539 = T84[1'h0:1'h0];
  assign T540 = T541 ? PArraySorted_3_7 : PArraySorted_2_7;
  assign T541 = T84[1'h0:1'h0];
  assign T542 = T84[1'h1:1'h1];
  assign T543 = T84[2'h2:2'h2];
  assign T544 = {T559, T545};
  assign T545 = T558 ? PArraySorted_4_8 : T546;
  assign T546 = T557 ? T555 : T547;
  assign T547 = T554 ? PArraySorted_1_8 : PArraySorted_0_8;
  assign T724 = reset ? 1'h0 : T548;
  assign T548 = T550 ? 1'h1 : T549;
  assign T549 = T593 ? 1'h0 : PArraySorted_0_8;
  assign T550 = T552 & T551;
  assign T551 = requestsBits[4'h8:4'h8];
  assign T552 = T593 & T553;
  assign T553 = io_requests_8_priorityLevel == 3'h0;
  assign T554 = T84[1'h0:1'h0];
  assign T555 = T556 ? PArraySorted_3_8 : PArraySorted_2_8;
  assign T556 = T84[1'h0:1'h0];
  assign T557 = T84[1'h1:1'h1];
  assign T558 = T84[2'h2:2'h2];
  assign T559 = T572 ? PArraySorted_4_9 : T560;
  assign T560 = T571 ? T569 : T561;
  assign T561 = T568 ? PArraySorted_1_9 : PArraySorted_0_9;
  assign T725 = reset ? 1'h0 : T562;
  assign T562 = T564 ? 1'h1 : T563;
  assign T563 = T593 ? 1'h0 : PArraySorted_0_9;
  assign T564 = T566 & T565;
  assign T565 = requestsBits[4'h9:4'h9];
  assign T566 = T593 & T567;
  assign T567 = io_requests_9_priorityLevel == 3'h0;
  assign T568 = T84[1'h0:1'h0];
  assign T569 = T570 ? PArraySorted_3_9 : PArraySorted_2_9;
  assign T570 = T84[1'h0:1'h0];
  assign T571 = T84[1'h1:1'h1];
  assign T572 = T84[2'h2:2'h2];
  assign T573 = T591 ? passSelectL1 : T574;
  assign T574 = passSelectL0[4'h9:1'h0];
  assign passSelectL0 = T575;
  assign T575 = T593 ? T576 : 11'h0;
  assign T576 = T582 + T577;
  assign T577 = {T581, T578};
  assign T578 = {T580, T579};
  assign T579 = nextGrant[4'h9:4'h9];
  assign T580 = nextGrant[4'h8:1'h0];
  assign T581 = 1'h0;
  assign T582 = {T585, T583};
  assign T583 = ~ T584;
  assign T584 = T64;
  assign T585 = 1'h0;
  assign passSelectL1 = T586;
  assign T586 = T593 ? T587 : 10'h0;
  assign T587 = T589 + T726;
  assign T726 = {9'h0, T588};
  assign T588 = 1'h1;
  assign T589 = ~ T590;
  assign T590 = T64;
  assign T591 = passSelectL0[4'ha:4'ha];
  assign T592 = winner != 10'h0;
  assign T593 = T59 & T594;
  assign T594 = T6 ^ 1'h1;
  assign T727 = winGrant[4'h9:4'h8];
  assign T728 = T653[3'h7:3'h4];
  assign T729 = T651[2'h3:2'h2];
  assign T730 = T729 != 2'h0;
  assign T731 = T728 != 4'h0;
  assign T732 = T727 != 2'h0;
  assign io_resource_valid = T595;
  assign T595 = T596 & io_resource_ready;
  assign T596 = T614 ? T612 : T597;
  assign T597 = T611 ? T605 : T598;
  assign T598 = T604 ? T602 : T599;
  assign T599 = T600 ? io_requests_1_grant : io_requests_0_grant;
  assign T600 = T601[1'h0:1'h0];
  assign T601 = io_chosen;
  assign T602 = T603 ? io_requests_3_grant : io_requests_2_grant;
  assign T603 = T601[1'h0:1'h0];
  assign T604 = T601[1'h1:1'h1];
  assign T605 = T610 ? T608 : T606;
  assign T606 = T607 ? io_requests_5_grant : io_requests_4_grant;
  assign T607 = T601[1'h0:1'h0];
  assign T608 = T609 ? io_requests_7_grant : io_requests_6_grant;
  assign T609 = T601[1'h0:1'h0];
  assign T610 = T601[1'h1:1'h1];
  assign T611 = T601[2'h2:2'h2];
  assign T612 = T613 ? io_requests_9_grant : io_requests_8_grant;
  assign T613 = T601[1'h0:1'h0];
  assign T614 = T601[2'h3:2'h3];
  assign io_requests_0_grant = T615;
  assign T615 = T616 & io_resource_ready;
  assign T616 = T617;
  assign T617 = winGrant[1'h0:1'h0];
  assign io_requests_1_grant = T618;
  assign T618 = T619 & io_resource_ready;
  assign T619 = T620;
  assign T620 = winGrant[1'h1:1'h1];
  assign io_requests_2_grant = T621;
  assign T621 = T622 & io_resource_ready;
  assign T622 = T623;
  assign T623 = winGrant[2'h2:2'h2];
  assign io_requests_3_grant = T624;
  assign T624 = T625 & io_resource_ready;
  assign T625 = T626;
  assign T626 = winGrant[2'h3:2'h3];
  assign io_requests_4_grant = T627;
  assign T627 = T628 & io_resource_ready;
  assign T628 = T629;
  assign T629 = winGrant[3'h4:3'h4];
  assign io_requests_5_grant = T630;
  assign T630 = T631 & io_resource_ready;
  assign T631 = T632;
  assign T632 = winGrant[3'h5:3'h5];
  assign io_requests_6_grant = T633;
  assign T633 = T634 & io_resource_ready;
  assign T634 = T635;
  assign T635 = winGrant[3'h6:3'h6];
  assign io_requests_7_grant = T636;
  assign T636 = T637 & io_resource_ready;
  assign T637 = T638;
  assign T638 = winGrant[3'h7:3'h7];
  assign io_requests_8_grant = T639;
  assign T639 = T640 & io_resource_ready;
  assign T640 = T641;
  assign T641 = winGrant[4'h8:4'h8];
  assign io_requests_9_grant = T642;
  assign T642 = T643 & io_resource_ready;
  assign T643 = T644;
  assign T644 = winGrant[4'h9:4'h9];

  always @(posedge clk) begin
    if(reset) begin
      nextGrant <= 10'h200;
    end else if(T593) begin
      nextGrant <= winGrant;
    end else if(T5) begin
      nextGrant <= winGrant;
    end
    if(reset) begin
      PArraySorted_0_0 <= 1'h0;
    end else if(T73) begin
      PArraySorted_0_0 <= 1'h1;
    end else if(T593) begin
      PArraySorted_0_0 <= 1'h0;
    end
    if(reset) begin
      PArraySorted_1_0 <= 1'h0;
    end else if(T79) begin
      PArraySorted_1_0 <= 1'h1;
    end else if(T593) begin
      PArraySorted_1_0 <= 1'h0;
    end
    if(reset) begin
      PArraySorted_1_1 <= 1'h0;
    end else if(T130) begin
      PArraySorted_1_1 <= 1'h1;
    end else if(T593) begin
      PArraySorted_1_1 <= 1'h0;
    end
    if(reset) begin
      PArraySorted_1_2 <= 1'h0;
    end else if(T138) begin
      PArraySorted_1_2 <= 1'h1;
    end else if(T593) begin
      PArraySorted_1_2 <= 1'h0;
    end
    if(reset) begin
      PArraySorted_1_3 <= 1'h0;
    end else if(T146) begin
      PArraySorted_1_3 <= 1'h1;
    end else if(T593) begin
      PArraySorted_1_3 <= 1'h0;
    end
    if(reset) begin
      PArraySorted_1_4 <= 1'h0;
    end else if(T154) begin
      PArraySorted_1_4 <= 1'h1;
    end else if(T593) begin
      PArraySorted_1_4 <= 1'h0;
    end
    if(reset) begin
      PArraySorted_1_5 <= 1'h0;
    end else if(T162) begin
      PArraySorted_1_5 <= 1'h1;
    end else if(T593) begin
      PArraySorted_1_5 <= 1'h0;
    end
    if(reset) begin
      PArraySorted_1_6 <= 1'h0;
    end else if(T170) begin
      PArraySorted_1_6 <= 1'h1;
    end else if(T593) begin
      PArraySorted_1_6 <= 1'h0;
    end
    if(reset) begin
      PArraySorted_1_7 <= 1'h0;
    end else if(T178) begin
      PArraySorted_1_7 <= 1'h1;
    end else if(T593) begin
      PArraySorted_1_7 <= 1'h0;
    end
    if(reset) begin
      PArraySorted_1_8 <= 1'h0;
    end else if(T186) begin
      PArraySorted_1_8 <= 1'h1;
    end else if(T593) begin
      PArraySorted_1_8 <= 1'h0;
    end
    if(reset) begin
      PArraySorted_1_9 <= 1'h0;
    end else if(T194) begin
      PArraySorted_1_9 <= 1'h1;
    end else if(T593) begin
      PArraySorted_1_9 <= 1'h0;
    end
    if(reset) begin
      PArraySorted_2_0 <= 1'h0;
    end else if(T202) begin
      PArraySorted_2_0 <= 1'h1;
    end else if(T593) begin
      PArraySorted_2_0 <= 1'h0;
    end
    if(reset) begin
      PArraySorted_2_1 <= 1'h0;
    end else if(T210) begin
      PArraySorted_2_1 <= 1'h1;
    end else if(T593) begin
      PArraySorted_2_1 <= 1'h0;
    end
    if(reset) begin
      PArraySorted_2_2 <= 1'h0;
    end else if(T218) begin
      PArraySorted_2_2 <= 1'h1;
    end else if(T593) begin
      PArraySorted_2_2 <= 1'h0;
    end
    if(reset) begin
      PArraySorted_2_3 <= 1'h0;
    end else if(T226) begin
      PArraySorted_2_3 <= 1'h1;
    end else if(T593) begin
      PArraySorted_2_3 <= 1'h0;
    end
    if(reset) begin
      PArraySorted_2_4 <= 1'h0;
    end else if(T234) begin
      PArraySorted_2_4 <= 1'h1;
    end else if(T593) begin
      PArraySorted_2_4 <= 1'h0;
    end
    if(reset) begin
      PArraySorted_2_5 <= 1'h0;
    end else if(T242) begin
      PArraySorted_2_5 <= 1'h1;
    end else if(T593) begin
      PArraySorted_2_5 <= 1'h0;
    end
    if(reset) begin
      PArraySorted_2_6 <= 1'h0;
    end else if(T250) begin
      PArraySorted_2_6 <= 1'h1;
    end else if(T593) begin
      PArraySorted_2_6 <= 1'h0;
    end
    if(reset) begin
      PArraySorted_2_7 <= 1'h0;
    end else if(T258) begin
      PArraySorted_2_7 <= 1'h1;
    end else if(T593) begin
      PArraySorted_2_7 <= 1'h0;
    end
    if(reset) begin
      PArraySorted_2_8 <= 1'h0;
    end else if(T266) begin
      PArraySorted_2_8 <= 1'h1;
    end else if(T593) begin
      PArraySorted_2_8 <= 1'h0;
    end
    if(reset) begin
      PArraySorted_2_9 <= 1'h0;
    end else if(T274) begin
      PArraySorted_2_9 <= 1'h1;
    end else if(T593) begin
      PArraySorted_2_9 <= 1'h0;
    end
    if(reset) begin
      PArraySorted_3_0 <= 1'h0;
    end else if(T282) begin
      PArraySorted_3_0 <= 1'h1;
    end else if(T593) begin
      PArraySorted_3_0 <= 1'h0;
    end
    if(reset) begin
      PArraySorted_3_1 <= 1'h0;
    end else if(T290) begin
      PArraySorted_3_1 <= 1'h1;
    end else if(T593) begin
      PArraySorted_3_1 <= 1'h0;
    end
    if(reset) begin
      PArraySorted_3_2 <= 1'h0;
    end else if(T298) begin
      PArraySorted_3_2 <= 1'h1;
    end else if(T593) begin
      PArraySorted_3_2 <= 1'h0;
    end
    if(reset) begin
      PArraySorted_3_3 <= 1'h0;
    end else if(T306) begin
      PArraySorted_3_3 <= 1'h1;
    end else if(T593) begin
      PArraySorted_3_3 <= 1'h0;
    end
    if(reset) begin
      PArraySorted_3_4 <= 1'h0;
    end else if(T314) begin
      PArraySorted_3_4 <= 1'h1;
    end else if(T593) begin
      PArraySorted_3_4 <= 1'h0;
    end
    if(reset) begin
      PArraySorted_3_5 <= 1'h0;
    end else if(T322) begin
      PArraySorted_3_5 <= 1'h1;
    end else if(T593) begin
      PArraySorted_3_5 <= 1'h0;
    end
    if(reset) begin
      PArraySorted_3_6 <= 1'h0;
    end else if(T330) begin
      PArraySorted_3_6 <= 1'h1;
    end else if(T593) begin
      PArraySorted_3_6 <= 1'h0;
    end
    if(reset) begin
      PArraySorted_3_7 <= 1'h0;
    end else if(T338) begin
      PArraySorted_3_7 <= 1'h1;
    end else if(T593) begin
      PArraySorted_3_7 <= 1'h0;
    end
    if(reset) begin
      PArraySorted_3_8 <= 1'h0;
    end else if(T346) begin
      PArraySorted_3_8 <= 1'h1;
    end else if(T593) begin
      PArraySorted_3_8 <= 1'h0;
    end
    if(reset) begin
      PArraySorted_3_9 <= 1'h0;
    end else if(T354) begin
      PArraySorted_3_9 <= 1'h1;
    end else if(T593) begin
      PArraySorted_3_9 <= 1'h0;
    end
    if(reset) begin
      PArraySorted_4_1 <= 1'h0;
    end else if(T364) begin
      PArraySorted_4_1 <= 1'h1;
    end else if(T593) begin
      PArraySorted_4_1 <= 1'h0;
    end
    if(reset) begin
      PArraySorted_4_2 <= 1'h0;
    end else if(T372) begin
      PArraySorted_4_2 <= 1'h1;
    end else if(T593) begin
      PArraySorted_4_2 <= 1'h0;
    end
    if(reset) begin
      PArraySorted_4_3 <= 1'h0;
    end else if(T380) begin
      PArraySorted_4_3 <= 1'h1;
    end else if(T593) begin
      PArraySorted_4_3 <= 1'h0;
    end
    if(reset) begin
      PArraySorted_4_4 <= 1'h0;
    end else if(T388) begin
      PArraySorted_4_4 <= 1'h1;
    end else if(T593) begin
      PArraySorted_4_4 <= 1'h0;
    end
    if(reset) begin
      PArraySorted_4_5 <= 1'h0;
    end else if(T396) begin
      PArraySorted_4_5 <= 1'h1;
    end else if(T593) begin
      PArraySorted_4_5 <= 1'h0;
    end
    if(reset) begin
      PArraySorted_4_6 <= 1'h0;
    end else if(T404) begin
      PArraySorted_4_6 <= 1'h1;
    end else if(T593) begin
      PArraySorted_4_6 <= 1'h0;
    end
    if(reset) begin
      PArraySorted_4_7 <= 1'h0;
    end else if(T412) begin
      PArraySorted_4_7 <= 1'h1;
    end else if(T593) begin
      PArraySorted_4_7 <= 1'h0;
    end
    if(reset) begin
      PArraySorted_4_8 <= 1'h0;
    end else if(T420) begin
      PArraySorted_4_8 <= 1'h1;
    end else if(T593) begin
      PArraySorted_4_8 <= 1'h0;
    end
    if(reset) begin
      PArraySorted_4_9 <= 1'h0;
    end else if(T428) begin
      PArraySorted_4_9 <= 1'h1;
    end else if(T593) begin
      PArraySorted_4_9 <= 1'h0;
    end
    if(reset) begin
      PArraySorted_4_0 <= 1'h0;
    end else if(T437) begin
      PArraySorted_4_0 <= 1'h1;
    end else if(T593) begin
      PArraySorted_4_0 <= 1'h0;
    end
    if(reset) begin
      PArraySorted_0_1 <= 1'h0;
    end else if(T447) begin
      PArraySorted_0_1 <= 1'h1;
    end else if(T593) begin
      PArraySorted_0_1 <= 1'h0;
    end
    if(reset) begin
      PArraySorted_0_2 <= 1'h0;
    end else if(T461) begin
      PArraySorted_0_2 <= 1'h1;
    end else if(T593) begin
      PArraySorted_0_2 <= 1'h0;
    end
    if(reset) begin
      PArraySorted_0_3 <= 1'h0;
    end else if(T476) begin
      PArraySorted_0_3 <= 1'h1;
    end else if(T593) begin
      PArraySorted_0_3 <= 1'h0;
    end
    if(reset) begin
      PArraySorted_0_4 <= 1'h0;
    end else if(T490) begin
      PArraySorted_0_4 <= 1'h1;
    end else if(T593) begin
      PArraySorted_0_4 <= 1'h0;
    end
    if(reset) begin
      PArraySorted_0_5 <= 1'h0;
    end else if(T507) begin
      PArraySorted_0_5 <= 1'h1;
    end else if(T593) begin
      PArraySorted_0_5 <= 1'h0;
    end
    if(reset) begin
      PArraySorted_0_6 <= 1'h0;
    end else if(T521) begin
      PArraySorted_0_6 <= 1'h1;
    end else if(T593) begin
      PArraySorted_0_6 <= 1'h0;
    end
    if(reset) begin
      PArraySorted_0_7 <= 1'h0;
    end else if(T535) begin
      PArraySorted_0_7 <= 1'h1;
    end else if(T593) begin
      PArraySorted_0_7 <= 1'h0;
    end
    if(reset) begin
      PArraySorted_0_8 <= 1'h0;
    end else if(T550) begin
      PArraySorted_0_8 <= 1'h1;
    end else if(T593) begin
      PArraySorted_0_8 <= 1'h0;
    end
    if(reset) begin
      PArraySorted_0_9 <= 1'h0;
    end else if(T564) begin
      PArraySorted_0_9 <= 1'h1;
    end else if(T593) begin
      PArraySorted_0_9 <= 1'h0;
    end
  end
endmodule

module SwitchAllocator_0(input clk, input reset,
    input  io_requests_4_9_releaseLock,
    output io_requests_4_9_grant,
    input  io_requests_4_9_request,
    input [2:0] io_requests_4_9_priorityLevel,
    input  io_requests_4_8_releaseLock,
    output io_requests_4_8_grant,
    input  io_requests_4_8_request,
    input [2:0] io_requests_4_8_priorityLevel,
    input  io_requests_4_7_releaseLock,
    output io_requests_4_7_grant,
    input  io_requests_4_7_request,
    input [2:0] io_requests_4_7_priorityLevel,
    input  io_requests_4_6_releaseLock,
    output io_requests_4_6_grant,
    input  io_requests_4_6_request,
    input [2:0] io_requests_4_6_priorityLevel,
    input  io_requests_4_5_releaseLock,
    output io_requests_4_5_grant,
    input  io_requests_4_5_request,
    input [2:0] io_requests_4_5_priorityLevel,
    input  io_requests_4_4_releaseLock,
    output io_requests_4_4_grant,
    input  io_requests_4_4_request,
    input [2:0] io_requests_4_4_priorityLevel,
    input  io_requests_4_3_releaseLock,
    output io_requests_4_3_grant,
    input  io_requests_4_3_request,
    input [2:0] io_requests_4_3_priorityLevel,
    input  io_requests_4_2_releaseLock,
    output io_requests_4_2_grant,
    input  io_requests_4_2_request,
    input [2:0] io_requests_4_2_priorityLevel,
    input  io_requests_4_1_releaseLock,
    output io_requests_4_1_grant,
    input  io_requests_4_1_request,
    input [2:0] io_requests_4_1_priorityLevel,
    input  io_requests_4_0_releaseLock,
    output io_requests_4_0_grant,
    input  io_requests_4_0_request,
    input [2:0] io_requests_4_0_priorityLevel,
    input  io_requests_3_9_releaseLock,
    output io_requests_3_9_grant,
    input  io_requests_3_9_request,
    input [2:0] io_requests_3_9_priorityLevel,
    input  io_requests_3_8_releaseLock,
    output io_requests_3_8_grant,
    input  io_requests_3_8_request,
    input [2:0] io_requests_3_8_priorityLevel,
    input  io_requests_3_7_releaseLock,
    output io_requests_3_7_grant,
    input  io_requests_3_7_request,
    input [2:0] io_requests_3_7_priorityLevel,
    input  io_requests_3_6_releaseLock,
    output io_requests_3_6_grant,
    input  io_requests_3_6_request,
    input [2:0] io_requests_3_6_priorityLevel,
    input  io_requests_3_5_releaseLock,
    output io_requests_3_5_grant,
    input  io_requests_3_5_request,
    input [2:0] io_requests_3_5_priorityLevel,
    input  io_requests_3_4_releaseLock,
    output io_requests_3_4_grant,
    input  io_requests_3_4_request,
    input [2:0] io_requests_3_4_priorityLevel,
    input  io_requests_3_3_releaseLock,
    output io_requests_3_3_grant,
    input  io_requests_3_3_request,
    input [2:0] io_requests_3_3_priorityLevel,
    input  io_requests_3_2_releaseLock,
    output io_requests_3_2_grant,
    input  io_requests_3_2_request,
    input [2:0] io_requests_3_2_priorityLevel,
    input  io_requests_3_1_releaseLock,
    output io_requests_3_1_grant,
    input  io_requests_3_1_request,
    input [2:0] io_requests_3_1_priorityLevel,
    input  io_requests_3_0_releaseLock,
    output io_requests_3_0_grant,
    input  io_requests_3_0_request,
    input [2:0] io_requests_3_0_priorityLevel,
    input  io_requests_2_9_releaseLock,
    output io_requests_2_9_grant,
    input  io_requests_2_9_request,
    input [2:0] io_requests_2_9_priorityLevel,
    input  io_requests_2_8_releaseLock,
    output io_requests_2_8_grant,
    input  io_requests_2_8_request,
    input [2:0] io_requests_2_8_priorityLevel,
    input  io_requests_2_7_releaseLock,
    output io_requests_2_7_grant,
    input  io_requests_2_7_request,
    input [2:0] io_requests_2_7_priorityLevel,
    input  io_requests_2_6_releaseLock,
    output io_requests_2_6_grant,
    input  io_requests_2_6_request,
    input [2:0] io_requests_2_6_priorityLevel,
    input  io_requests_2_5_releaseLock,
    output io_requests_2_5_grant,
    input  io_requests_2_5_request,
    input [2:0] io_requests_2_5_priorityLevel,
    input  io_requests_2_4_releaseLock,
    output io_requests_2_4_grant,
    input  io_requests_2_4_request,
    input [2:0] io_requests_2_4_priorityLevel,
    input  io_requests_2_3_releaseLock,
    output io_requests_2_3_grant,
    input  io_requests_2_3_request,
    input [2:0] io_requests_2_3_priorityLevel,
    input  io_requests_2_2_releaseLock,
    output io_requests_2_2_grant,
    input  io_requests_2_2_request,
    input [2:0] io_requests_2_2_priorityLevel,
    input  io_requests_2_1_releaseLock,
    output io_requests_2_1_grant,
    input  io_requests_2_1_request,
    input [2:0] io_requests_2_1_priorityLevel,
    input  io_requests_2_0_releaseLock,
    output io_requests_2_0_grant,
    input  io_requests_2_0_request,
    input [2:0] io_requests_2_0_priorityLevel,
    input  io_requests_1_9_releaseLock,
    output io_requests_1_9_grant,
    input  io_requests_1_9_request,
    input [2:0] io_requests_1_9_priorityLevel,
    input  io_requests_1_8_releaseLock,
    output io_requests_1_8_grant,
    input  io_requests_1_8_request,
    input [2:0] io_requests_1_8_priorityLevel,
    input  io_requests_1_7_releaseLock,
    output io_requests_1_7_grant,
    input  io_requests_1_7_request,
    input [2:0] io_requests_1_7_priorityLevel,
    input  io_requests_1_6_releaseLock,
    output io_requests_1_6_grant,
    input  io_requests_1_6_request,
    input [2:0] io_requests_1_6_priorityLevel,
    input  io_requests_1_5_releaseLock,
    output io_requests_1_5_grant,
    input  io_requests_1_5_request,
    input [2:0] io_requests_1_5_priorityLevel,
    input  io_requests_1_4_releaseLock,
    output io_requests_1_4_grant,
    input  io_requests_1_4_request,
    input [2:0] io_requests_1_4_priorityLevel,
    input  io_requests_1_3_releaseLock,
    output io_requests_1_3_grant,
    input  io_requests_1_3_request,
    input [2:0] io_requests_1_3_priorityLevel,
    input  io_requests_1_2_releaseLock,
    output io_requests_1_2_grant,
    input  io_requests_1_2_request,
    input [2:0] io_requests_1_2_priorityLevel,
    input  io_requests_1_1_releaseLock,
    output io_requests_1_1_grant,
    input  io_requests_1_1_request,
    input [2:0] io_requests_1_1_priorityLevel,
    input  io_requests_1_0_releaseLock,
    output io_requests_1_0_grant,
    input  io_requests_1_0_request,
    input [2:0] io_requests_1_0_priorityLevel,
    input  io_requests_0_9_releaseLock,
    output io_requests_0_9_grant,
    input  io_requests_0_9_request,
    input [2:0] io_requests_0_9_priorityLevel,
    input  io_requests_0_8_releaseLock,
    output io_requests_0_8_grant,
    input  io_requests_0_8_request,
    input [2:0] io_requests_0_8_priorityLevel,
    input  io_requests_0_7_releaseLock,
    output io_requests_0_7_grant,
    input  io_requests_0_7_request,
    input [2:0] io_requests_0_7_priorityLevel,
    input  io_requests_0_6_releaseLock,
    output io_requests_0_6_grant,
    input  io_requests_0_6_request,
    input [2:0] io_requests_0_6_priorityLevel,
    input  io_requests_0_5_releaseLock,
    output io_requests_0_5_grant,
    input  io_requests_0_5_request,
    input [2:0] io_requests_0_5_priorityLevel,
    input  io_requests_0_4_releaseLock,
    output io_requests_0_4_grant,
    input  io_requests_0_4_request,
    input [2:0] io_requests_0_4_priorityLevel,
    input  io_requests_0_3_releaseLock,
    output io_requests_0_3_grant,
    input  io_requests_0_3_request,
    input [2:0] io_requests_0_3_priorityLevel,
    input  io_requests_0_2_releaseLock,
    output io_requests_0_2_grant,
    input  io_requests_0_2_request,
    input [2:0] io_requests_0_2_priorityLevel,
    input  io_requests_0_1_releaseLock,
    output io_requests_0_1_grant,
    input  io_requests_0_1_request,
    input [2:0] io_requests_0_1_priorityLevel,
    input  io_requests_0_0_releaseLock,
    output io_requests_0_0_grant,
    input  io_requests_0_0_request,
    input [2:0] io_requests_0_0_priorityLevel,
    input  io_resources_4_ready,
    output io_resources_4_valid,
    input  io_resources_3_ready,
    output io_resources_3_valid,
    input  io_resources_2_ready,
    output io_resources_2_valid,
    input  io_resources_1_ready,
    output io_resources_1_valid,
    input  io_resources_0_ready,
    output io_resources_0_valid,
    output[3:0] io_chosens_4,
    output[3:0] io_chosens_3,
    output[3:0] io_chosens_2,
    output[3:0] io_chosens_1,
    output[3:0] io_chosens_0
);

  wire RRArbiterPriority_io_requests_9_grant;
  wire RRArbiterPriority_io_requests_8_grant;
  wire RRArbiterPriority_io_requests_7_grant;
  wire RRArbiterPriority_io_requests_6_grant;
  wire RRArbiterPriority_io_requests_5_grant;
  wire RRArbiterPriority_io_requests_4_grant;
  wire RRArbiterPriority_io_requests_3_grant;
  wire RRArbiterPriority_io_requests_2_grant;
  wire RRArbiterPriority_io_requests_1_grant;
  wire RRArbiterPriority_io_requests_0_grant;
  wire RRArbiterPriority_io_resource_valid;
  wire[3:0] RRArbiterPriority_io_chosen;
  wire RRArbiterPriority_1_io_requests_9_grant;
  wire RRArbiterPriority_1_io_requests_8_grant;
  wire RRArbiterPriority_1_io_requests_7_grant;
  wire RRArbiterPriority_1_io_requests_6_grant;
  wire RRArbiterPriority_1_io_requests_5_grant;
  wire RRArbiterPriority_1_io_requests_4_grant;
  wire RRArbiterPriority_1_io_requests_3_grant;
  wire RRArbiterPriority_1_io_requests_2_grant;
  wire RRArbiterPriority_1_io_requests_1_grant;
  wire RRArbiterPriority_1_io_requests_0_grant;
  wire RRArbiterPriority_1_io_resource_valid;
  wire[3:0] RRArbiterPriority_1_io_chosen;
  wire RRArbiterPriority_2_io_requests_9_grant;
  wire RRArbiterPriority_2_io_requests_8_grant;
  wire RRArbiterPriority_2_io_requests_7_grant;
  wire RRArbiterPriority_2_io_requests_6_grant;
  wire RRArbiterPriority_2_io_requests_5_grant;
  wire RRArbiterPriority_2_io_requests_4_grant;
  wire RRArbiterPriority_2_io_requests_3_grant;
  wire RRArbiterPriority_2_io_requests_2_grant;
  wire RRArbiterPriority_2_io_requests_1_grant;
  wire RRArbiterPriority_2_io_requests_0_grant;
  wire RRArbiterPriority_2_io_resource_valid;
  wire[3:0] RRArbiterPriority_2_io_chosen;
  wire RRArbiterPriority_3_io_requests_9_grant;
  wire RRArbiterPriority_3_io_requests_8_grant;
  wire RRArbiterPriority_3_io_requests_7_grant;
  wire RRArbiterPriority_3_io_requests_6_grant;
  wire RRArbiterPriority_3_io_requests_5_grant;
  wire RRArbiterPriority_3_io_requests_4_grant;
  wire RRArbiterPriority_3_io_requests_3_grant;
  wire RRArbiterPriority_3_io_requests_2_grant;
  wire RRArbiterPriority_3_io_requests_1_grant;
  wire RRArbiterPriority_3_io_requests_0_grant;
  wire RRArbiterPriority_3_io_resource_valid;
  wire[3:0] RRArbiterPriority_3_io_chosen;
  wire RRArbiterPriority_4_io_requests_9_grant;
  wire RRArbiterPriority_4_io_requests_8_grant;
  wire RRArbiterPriority_4_io_requests_7_grant;
  wire RRArbiterPriority_4_io_requests_6_grant;
  wire RRArbiterPriority_4_io_requests_5_grant;
  wire RRArbiterPriority_4_io_requests_4_grant;
  wire RRArbiterPriority_4_io_requests_3_grant;
  wire RRArbiterPriority_4_io_requests_2_grant;
  wire RRArbiterPriority_4_io_requests_1_grant;
  wire RRArbiterPriority_4_io_requests_0_grant;
  wire RRArbiterPriority_4_io_resource_valid;
  wire[3:0] RRArbiterPriority_4_io_chosen;


  assign io_chosens_0 = RRArbiterPriority_io_chosen;
  assign io_chosens_1 = RRArbiterPriority_1_io_chosen;
  assign io_chosens_2 = RRArbiterPriority_2_io_chosen;
  assign io_chosens_3 = RRArbiterPriority_3_io_chosen;
  assign io_chosens_4 = RRArbiterPriority_4_io_chosen;
  assign io_resources_0_valid = RRArbiterPriority_io_resource_valid;
  assign io_resources_1_valid = RRArbiterPriority_1_io_resource_valid;
  assign io_resources_2_valid = RRArbiterPriority_2_io_resource_valid;
  assign io_resources_3_valid = RRArbiterPriority_3_io_resource_valid;
  assign io_resources_4_valid = RRArbiterPriority_4_io_resource_valid;
  assign io_requests_0_0_grant = RRArbiterPriority_io_requests_0_grant;
  assign io_requests_0_1_grant = RRArbiterPriority_io_requests_1_grant;
  assign io_requests_0_2_grant = RRArbiterPriority_io_requests_2_grant;
  assign io_requests_0_3_grant = RRArbiterPriority_io_requests_3_grant;
  assign io_requests_0_4_grant = RRArbiterPriority_io_requests_4_grant;
  assign io_requests_0_5_grant = RRArbiterPriority_io_requests_5_grant;
  assign io_requests_0_6_grant = RRArbiterPriority_io_requests_6_grant;
  assign io_requests_0_7_grant = RRArbiterPriority_io_requests_7_grant;
  assign io_requests_0_8_grant = RRArbiterPriority_io_requests_8_grant;
  assign io_requests_0_9_grant = RRArbiterPriority_io_requests_9_grant;
  assign io_requests_1_0_grant = RRArbiterPriority_1_io_requests_0_grant;
  assign io_requests_1_1_grant = RRArbiterPriority_1_io_requests_1_grant;
  assign io_requests_1_2_grant = RRArbiterPriority_1_io_requests_2_grant;
  assign io_requests_1_3_grant = RRArbiterPriority_1_io_requests_3_grant;
  assign io_requests_1_4_grant = RRArbiterPriority_1_io_requests_4_grant;
  assign io_requests_1_5_grant = RRArbiterPriority_1_io_requests_5_grant;
  assign io_requests_1_6_grant = RRArbiterPriority_1_io_requests_6_grant;
  assign io_requests_1_7_grant = RRArbiterPriority_1_io_requests_7_grant;
  assign io_requests_1_8_grant = RRArbiterPriority_1_io_requests_8_grant;
  assign io_requests_1_9_grant = RRArbiterPriority_1_io_requests_9_grant;
  assign io_requests_2_0_grant = RRArbiterPriority_2_io_requests_0_grant;
  assign io_requests_2_1_grant = RRArbiterPriority_2_io_requests_1_grant;
  assign io_requests_2_2_grant = RRArbiterPriority_2_io_requests_2_grant;
  assign io_requests_2_3_grant = RRArbiterPriority_2_io_requests_3_grant;
  assign io_requests_2_4_grant = RRArbiterPriority_2_io_requests_4_grant;
  assign io_requests_2_5_grant = RRArbiterPriority_2_io_requests_5_grant;
  assign io_requests_2_6_grant = RRArbiterPriority_2_io_requests_6_grant;
  assign io_requests_2_7_grant = RRArbiterPriority_2_io_requests_7_grant;
  assign io_requests_2_8_grant = RRArbiterPriority_2_io_requests_8_grant;
  assign io_requests_2_9_grant = RRArbiterPriority_2_io_requests_9_grant;
  assign io_requests_3_0_grant = RRArbiterPriority_3_io_requests_0_grant;
  assign io_requests_3_1_grant = RRArbiterPriority_3_io_requests_1_grant;
  assign io_requests_3_2_grant = RRArbiterPriority_3_io_requests_2_grant;
  assign io_requests_3_3_grant = RRArbiterPriority_3_io_requests_3_grant;
  assign io_requests_3_4_grant = RRArbiterPriority_3_io_requests_4_grant;
  assign io_requests_3_5_grant = RRArbiterPriority_3_io_requests_5_grant;
  assign io_requests_3_6_grant = RRArbiterPriority_3_io_requests_6_grant;
  assign io_requests_3_7_grant = RRArbiterPriority_3_io_requests_7_grant;
  assign io_requests_3_8_grant = RRArbiterPriority_3_io_requests_8_grant;
  assign io_requests_3_9_grant = RRArbiterPriority_3_io_requests_9_grant;
  assign io_requests_4_0_grant = RRArbiterPriority_4_io_requests_0_grant;
  assign io_requests_4_1_grant = RRArbiterPriority_4_io_requests_1_grant;
  assign io_requests_4_2_grant = RRArbiterPriority_4_io_requests_2_grant;
  assign io_requests_4_3_grant = RRArbiterPriority_4_io_requests_3_grant;
  assign io_requests_4_4_grant = RRArbiterPriority_4_io_requests_4_grant;
  assign io_requests_4_5_grant = RRArbiterPriority_4_io_requests_5_grant;
  assign io_requests_4_6_grant = RRArbiterPriority_4_io_requests_6_grant;
  assign io_requests_4_7_grant = RRArbiterPriority_4_io_requests_7_grant;
  assign io_requests_4_8_grant = RRArbiterPriority_4_io_requests_8_grant;
  assign io_requests_4_9_grant = RRArbiterPriority_4_io_requests_9_grant;
  RRArbiterPriority RRArbiterPriority(.clk(clk), .reset(reset),
       .io_requests_9_releaseLock( io_requests_0_9_releaseLock ),
       .io_requests_9_grant( RRArbiterPriority_io_requests_9_grant ),
       .io_requests_9_request( io_requests_0_9_request ),
       .io_requests_9_priorityLevel( io_requests_0_9_priorityLevel ),
       .io_requests_8_releaseLock( io_requests_0_8_releaseLock ),
       .io_requests_8_grant( RRArbiterPriority_io_requests_8_grant ),
       .io_requests_8_request( io_requests_0_8_request ),
       .io_requests_8_priorityLevel( io_requests_0_8_priorityLevel ),
       .io_requests_7_releaseLock( io_requests_0_7_releaseLock ),
       .io_requests_7_grant( RRArbiterPriority_io_requests_7_grant ),
       .io_requests_7_request( io_requests_0_7_request ),
       .io_requests_7_priorityLevel( io_requests_0_7_priorityLevel ),
       .io_requests_6_releaseLock( io_requests_0_6_releaseLock ),
       .io_requests_6_grant( RRArbiterPriority_io_requests_6_grant ),
       .io_requests_6_request( io_requests_0_6_request ),
       .io_requests_6_priorityLevel( io_requests_0_6_priorityLevel ),
       .io_requests_5_releaseLock( io_requests_0_5_releaseLock ),
       .io_requests_5_grant( RRArbiterPriority_io_requests_5_grant ),
       .io_requests_5_request( io_requests_0_5_request ),
       .io_requests_5_priorityLevel( io_requests_0_5_priorityLevel ),
       .io_requests_4_releaseLock( io_requests_0_4_releaseLock ),
       .io_requests_4_grant( RRArbiterPriority_io_requests_4_grant ),
       .io_requests_4_request( io_requests_0_4_request ),
       .io_requests_4_priorityLevel( io_requests_0_4_priorityLevel ),
       .io_requests_3_releaseLock( io_requests_0_3_releaseLock ),
       .io_requests_3_grant( RRArbiterPriority_io_requests_3_grant ),
       .io_requests_3_request( io_requests_0_3_request ),
       .io_requests_3_priorityLevel( io_requests_0_3_priorityLevel ),
       .io_requests_2_releaseLock( io_requests_0_2_releaseLock ),
       .io_requests_2_grant( RRArbiterPriority_io_requests_2_grant ),
       .io_requests_2_request( io_requests_0_2_request ),
       .io_requests_2_priorityLevel( io_requests_0_2_priorityLevel ),
       .io_requests_1_releaseLock( io_requests_0_1_releaseLock ),
       .io_requests_1_grant( RRArbiterPriority_io_requests_1_grant ),
       .io_requests_1_request( io_requests_0_1_request ),
       .io_requests_1_priorityLevel( io_requests_0_1_priorityLevel ),
       .io_requests_0_releaseLock( io_requests_0_0_releaseLock ),
       .io_requests_0_grant( RRArbiterPriority_io_requests_0_grant ),
       .io_requests_0_request( io_requests_0_0_request ),
       .io_requests_0_priorityLevel( io_requests_0_0_priorityLevel ),
       .io_resource_ready( io_resources_0_ready ),
       .io_resource_valid( RRArbiterPriority_io_resource_valid ),
       .io_chosen( RRArbiterPriority_io_chosen )
  );
  RRArbiterPriority RRArbiterPriority_1(.clk(clk), .reset(reset),
       .io_requests_9_releaseLock( io_requests_1_9_releaseLock ),
       .io_requests_9_grant( RRArbiterPriority_1_io_requests_9_grant ),
       .io_requests_9_request( io_requests_1_9_request ),
       .io_requests_9_priorityLevel( io_requests_1_9_priorityLevel ),
       .io_requests_8_releaseLock( io_requests_1_8_releaseLock ),
       .io_requests_8_grant( RRArbiterPriority_1_io_requests_8_grant ),
       .io_requests_8_request( io_requests_1_8_request ),
       .io_requests_8_priorityLevel( io_requests_1_8_priorityLevel ),
       .io_requests_7_releaseLock( io_requests_1_7_releaseLock ),
       .io_requests_7_grant( RRArbiterPriority_1_io_requests_7_grant ),
       .io_requests_7_request( io_requests_1_7_request ),
       .io_requests_7_priorityLevel( io_requests_1_7_priorityLevel ),
       .io_requests_6_releaseLock( io_requests_1_6_releaseLock ),
       .io_requests_6_grant( RRArbiterPriority_1_io_requests_6_grant ),
       .io_requests_6_request( io_requests_1_6_request ),
       .io_requests_6_priorityLevel( io_requests_1_6_priorityLevel ),
       .io_requests_5_releaseLock( io_requests_1_5_releaseLock ),
       .io_requests_5_grant( RRArbiterPriority_1_io_requests_5_grant ),
       .io_requests_5_request( io_requests_1_5_request ),
       .io_requests_5_priorityLevel( io_requests_1_5_priorityLevel ),
       .io_requests_4_releaseLock( io_requests_1_4_releaseLock ),
       .io_requests_4_grant( RRArbiterPriority_1_io_requests_4_grant ),
       .io_requests_4_request( io_requests_1_4_request ),
       .io_requests_4_priorityLevel( io_requests_1_4_priorityLevel ),
       .io_requests_3_releaseLock( io_requests_1_3_releaseLock ),
       .io_requests_3_grant( RRArbiterPriority_1_io_requests_3_grant ),
       .io_requests_3_request( io_requests_1_3_request ),
       .io_requests_3_priorityLevel( io_requests_1_3_priorityLevel ),
       .io_requests_2_releaseLock( io_requests_1_2_releaseLock ),
       .io_requests_2_grant( RRArbiterPriority_1_io_requests_2_grant ),
       .io_requests_2_request( io_requests_1_2_request ),
       .io_requests_2_priorityLevel( io_requests_1_2_priorityLevel ),
       .io_requests_1_releaseLock( io_requests_1_1_releaseLock ),
       .io_requests_1_grant( RRArbiterPriority_1_io_requests_1_grant ),
       .io_requests_1_request( io_requests_1_1_request ),
       .io_requests_1_priorityLevel( io_requests_1_1_priorityLevel ),
       .io_requests_0_releaseLock( io_requests_1_0_releaseLock ),
       .io_requests_0_grant( RRArbiterPriority_1_io_requests_0_grant ),
       .io_requests_0_request( io_requests_1_0_request ),
       .io_requests_0_priorityLevel( io_requests_1_0_priorityLevel ),
       .io_resource_ready( io_resources_1_ready ),
       .io_resource_valid( RRArbiterPriority_1_io_resource_valid ),
       .io_chosen( RRArbiterPriority_1_io_chosen )
  );
  RRArbiterPriority RRArbiterPriority_2(.clk(clk), .reset(reset),
       .io_requests_9_releaseLock( io_requests_2_9_releaseLock ),
       .io_requests_9_grant( RRArbiterPriority_2_io_requests_9_grant ),
       .io_requests_9_request( io_requests_2_9_request ),
       .io_requests_9_priorityLevel( io_requests_2_9_priorityLevel ),
       .io_requests_8_releaseLock( io_requests_2_8_releaseLock ),
       .io_requests_8_grant( RRArbiterPriority_2_io_requests_8_grant ),
       .io_requests_8_request( io_requests_2_8_request ),
       .io_requests_8_priorityLevel( io_requests_2_8_priorityLevel ),
       .io_requests_7_releaseLock( io_requests_2_7_releaseLock ),
       .io_requests_7_grant( RRArbiterPriority_2_io_requests_7_grant ),
       .io_requests_7_request( io_requests_2_7_request ),
       .io_requests_7_priorityLevel( io_requests_2_7_priorityLevel ),
       .io_requests_6_releaseLock( io_requests_2_6_releaseLock ),
       .io_requests_6_grant( RRArbiterPriority_2_io_requests_6_grant ),
       .io_requests_6_request( io_requests_2_6_request ),
       .io_requests_6_priorityLevel( io_requests_2_6_priorityLevel ),
       .io_requests_5_releaseLock( io_requests_2_5_releaseLock ),
       .io_requests_5_grant( RRArbiterPriority_2_io_requests_5_grant ),
       .io_requests_5_request( io_requests_2_5_request ),
       .io_requests_5_priorityLevel( io_requests_2_5_priorityLevel ),
       .io_requests_4_releaseLock( io_requests_2_4_releaseLock ),
       .io_requests_4_grant( RRArbiterPriority_2_io_requests_4_grant ),
       .io_requests_4_request( io_requests_2_4_request ),
       .io_requests_4_priorityLevel( io_requests_2_4_priorityLevel ),
       .io_requests_3_releaseLock( io_requests_2_3_releaseLock ),
       .io_requests_3_grant( RRArbiterPriority_2_io_requests_3_grant ),
       .io_requests_3_request( io_requests_2_3_request ),
       .io_requests_3_priorityLevel( io_requests_2_3_priorityLevel ),
       .io_requests_2_releaseLock( io_requests_2_2_releaseLock ),
       .io_requests_2_grant( RRArbiterPriority_2_io_requests_2_grant ),
       .io_requests_2_request( io_requests_2_2_request ),
       .io_requests_2_priorityLevel( io_requests_2_2_priorityLevel ),
       .io_requests_1_releaseLock( io_requests_2_1_releaseLock ),
       .io_requests_1_grant( RRArbiterPriority_2_io_requests_1_grant ),
       .io_requests_1_request( io_requests_2_1_request ),
       .io_requests_1_priorityLevel( io_requests_2_1_priorityLevel ),
       .io_requests_0_releaseLock( io_requests_2_0_releaseLock ),
       .io_requests_0_grant( RRArbiterPriority_2_io_requests_0_grant ),
       .io_requests_0_request( io_requests_2_0_request ),
       .io_requests_0_priorityLevel( io_requests_2_0_priorityLevel ),
       .io_resource_ready( io_resources_2_ready ),
       .io_resource_valid( RRArbiterPriority_2_io_resource_valid ),
       .io_chosen( RRArbiterPriority_2_io_chosen )
  );
  RRArbiterPriority RRArbiterPriority_3(.clk(clk), .reset(reset),
       .io_requests_9_releaseLock( io_requests_3_9_releaseLock ),
       .io_requests_9_grant( RRArbiterPriority_3_io_requests_9_grant ),
       .io_requests_9_request( io_requests_3_9_request ),
       .io_requests_9_priorityLevel( io_requests_3_9_priorityLevel ),
       .io_requests_8_releaseLock( io_requests_3_8_releaseLock ),
       .io_requests_8_grant( RRArbiterPriority_3_io_requests_8_grant ),
       .io_requests_8_request( io_requests_3_8_request ),
       .io_requests_8_priorityLevel( io_requests_3_8_priorityLevel ),
       .io_requests_7_releaseLock( io_requests_3_7_releaseLock ),
       .io_requests_7_grant( RRArbiterPriority_3_io_requests_7_grant ),
       .io_requests_7_request( io_requests_3_7_request ),
       .io_requests_7_priorityLevel( io_requests_3_7_priorityLevel ),
       .io_requests_6_releaseLock( io_requests_3_6_releaseLock ),
       .io_requests_6_grant( RRArbiterPriority_3_io_requests_6_grant ),
       .io_requests_6_request( io_requests_3_6_request ),
       .io_requests_6_priorityLevel( io_requests_3_6_priorityLevel ),
       .io_requests_5_releaseLock( io_requests_3_5_releaseLock ),
       .io_requests_5_grant( RRArbiterPriority_3_io_requests_5_grant ),
       .io_requests_5_request( io_requests_3_5_request ),
       .io_requests_5_priorityLevel( io_requests_3_5_priorityLevel ),
       .io_requests_4_releaseLock( io_requests_3_4_releaseLock ),
       .io_requests_4_grant( RRArbiterPriority_3_io_requests_4_grant ),
       .io_requests_4_request( io_requests_3_4_request ),
       .io_requests_4_priorityLevel( io_requests_3_4_priorityLevel ),
       .io_requests_3_releaseLock( io_requests_3_3_releaseLock ),
       .io_requests_3_grant( RRArbiterPriority_3_io_requests_3_grant ),
       .io_requests_3_request( io_requests_3_3_request ),
       .io_requests_3_priorityLevel( io_requests_3_3_priorityLevel ),
       .io_requests_2_releaseLock( io_requests_3_2_releaseLock ),
       .io_requests_2_grant( RRArbiterPriority_3_io_requests_2_grant ),
       .io_requests_2_request( io_requests_3_2_request ),
       .io_requests_2_priorityLevel( io_requests_3_2_priorityLevel ),
       .io_requests_1_releaseLock( io_requests_3_1_releaseLock ),
       .io_requests_1_grant( RRArbiterPriority_3_io_requests_1_grant ),
       .io_requests_1_request( io_requests_3_1_request ),
       .io_requests_1_priorityLevel( io_requests_3_1_priorityLevel ),
       .io_requests_0_releaseLock( io_requests_3_0_releaseLock ),
       .io_requests_0_grant( RRArbiterPriority_3_io_requests_0_grant ),
       .io_requests_0_request( io_requests_3_0_request ),
       .io_requests_0_priorityLevel( io_requests_3_0_priorityLevel ),
       .io_resource_ready( io_resources_3_ready ),
       .io_resource_valid( RRArbiterPriority_3_io_resource_valid ),
       .io_chosen( RRArbiterPriority_3_io_chosen )
  );
  RRArbiterPriority RRArbiterPriority_4(.clk(clk), .reset(reset),
       .io_requests_9_releaseLock( io_requests_4_9_releaseLock ),
       .io_requests_9_grant( RRArbiterPriority_4_io_requests_9_grant ),
       .io_requests_9_request( io_requests_4_9_request ),
       .io_requests_9_priorityLevel( io_requests_4_9_priorityLevel ),
       .io_requests_8_releaseLock( io_requests_4_8_releaseLock ),
       .io_requests_8_grant( RRArbiterPriority_4_io_requests_8_grant ),
       .io_requests_8_request( io_requests_4_8_request ),
       .io_requests_8_priorityLevel( io_requests_4_8_priorityLevel ),
       .io_requests_7_releaseLock( io_requests_4_7_releaseLock ),
       .io_requests_7_grant( RRArbiterPriority_4_io_requests_7_grant ),
       .io_requests_7_request( io_requests_4_7_request ),
       .io_requests_7_priorityLevel( io_requests_4_7_priorityLevel ),
       .io_requests_6_releaseLock( io_requests_4_6_releaseLock ),
       .io_requests_6_grant( RRArbiterPriority_4_io_requests_6_grant ),
       .io_requests_6_request( io_requests_4_6_request ),
       .io_requests_6_priorityLevel( io_requests_4_6_priorityLevel ),
       .io_requests_5_releaseLock( io_requests_4_5_releaseLock ),
       .io_requests_5_grant( RRArbiterPriority_4_io_requests_5_grant ),
       .io_requests_5_request( io_requests_4_5_request ),
       .io_requests_5_priorityLevel( io_requests_4_5_priorityLevel ),
       .io_requests_4_releaseLock( io_requests_4_4_releaseLock ),
       .io_requests_4_grant( RRArbiterPriority_4_io_requests_4_grant ),
       .io_requests_4_request( io_requests_4_4_request ),
       .io_requests_4_priorityLevel( io_requests_4_4_priorityLevel ),
       .io_requests_3_releaseLock( io_requests_4_3_releaseLock ),
       .io_requests_3_grant( RRArbiterPriority_4_io_requests_3_grant ),
       .io_requests_3_request( io_requests_4_3_request ),
       .io_requests_3_priorityLevel( io_requests_4_3_priorityLevel ),
       .io_requests_2_releaseLock( io_requests_4_2_releaseLock ),
       .io_requests_2_grant( RRArbiterPriority_4_io_requests_2_grant ),
       .io_requests_2_request( io_requests_4_2_request ),
       .io_requests_2_priorityLevel( io_requests_4_2_priorityLevel ),
       .io_requests_1_releaseLock( io_requests_4_1_releaseLock ),
       .io_requests_1_grant( RRArbiterPriority_4_io_requests_1_grant ),
       .io_requests_1_request( io_requests_4_1_request ),
       .io_requests_1_priorityLevel( io_requests_4_1_priorityLevel ),
       .io_requests_0_releaseLock( io_requests_4_0_releaseLock ),
       .io_requests_0_grant( RRArbiterPriority_4_io_requests_0_grant ),
       .io_requests_0_request( io_requests_4_0_request ),
       .io_requests_0_priorityLevel( io_requests_4_0_priorityLevel ),
       .io_resource_ready( io_resources_4_ready ),
       .io_resource_valid( RRArbiterPriority_4_io_resource_valid ),
       .io_chosen( RRArbiterPriority_4_io_chosen )
  );
endmodule

module RRArbiter_1(input clk, input reset,
    input  io_requests_9_releaseLock,
    output io_requests_9_grant,
    input  io_requests_9_request,
    input [2:0] io_requests_9_priorityLevel,
    input  io_requests_8_releaseLock,
    output io_requests_8_grant,
    input  io_requests_8_request,
    input [2:0] io_requests_8_priorityLevel,
    input  io_requests_7_releaseLock,
    output io_requests_7_grant,
    input  io_requests_7_request,
    input [2:0] io_requests_7_priorityLevel,
    input  io_requests_6_releaseLock,
    output io_requests_6_grant,
    input  io_requests_6_request,
    input [2:0] io_requests_6_priorityLevel,
    input  io_requests_5_releaseLock,
    output io_requests_5_grant,
    input  io_requests_5_request,
    input [2:0] io_requests_5_priorityLevel,
    input  io_requests_4_releaseLock,
    output io_requests_4_grant,
    input  io_requests_4_request,
    input [2:0] io_requests_4_priorityLevel,
    input  io_requests_3_releaseLock,
    output io_requests_3_grant,
    input  io_requests_3_request,
    input [2:0] io_requests_3_priorityLevel,
    input  io_requests_2_releaseLock,
    output io_requests_2_grant,
    input  io_requests_2_request,
    input [2:0] io_requests_2_priorityLevel,
    input  io_requests_1_releaseLock,
    output io_requests_1_grant,
    input  io_requests_1_request,
    input [2:0] io_requests_1_priorityLevel,
    input  io_requests_0_releaseLock,
    output io_requests_0_grant,
    input  io_requests_0_request,
    input [2:0] io_requests_0_priorityLevel,
    input  io_resource_ready,
    output io_resource_valid,
    output[3:0] io_chosen
);

  wire[3:0] T127;
  wire[2:0] T128;
  wire[1:0] T129;
  wire T130;
  wire[1:0] T131;
  wire[1:0] T132;
  wire[3:0] T133;
  wire[3:0] T134;
  wire[7:0] T135;
  wire[7:0] T136;
  wire[9:0] winner;
  wire[9:0] T1;
  reg [9:0] nextGrant;
  wire[9:0] T137;
  wire[9:0] T2;
  wire[9:0] T3;
  wire T4;
  wire[9:0] T5;
  wire[9:0] requestsBits;
  wire[4:0] T6;
  wire[2:0] T7;
  wire[1:0] T8;
  wire T9;
  wire T10;
  wire T11;
  wire[1:0] T12;
  wire T13;
  wire T14;
  wire[4:0] T15;
  wire[2:0] T16;
  wire[1:0] T17;
  wire T18;
  wire T19;
  wire T20;
  wire[1:0] T21;
  wire T22;
  wire T23;
  wire[9:0] T24;
  wire[9:0] T25;
  wire[10:0] passSelectL0;
  wire[10:0] T26;
  wire[10:0] T27;
  wire[10:0] T28;
  wire[9:0] T29;
  wire T30;
  wire[8:0] T31;
  wire T32;
  wire[10:0] T33;
  wire[9:0] T34;
  wire T35;
  wire[9:0] passSelectL1;
  wire[9:0] T36;
  wire[9:0] T37;
  wire[9:0] T138;
  wire T38;
  wire[9:0] T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire lockRelease;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire[3:0] T49;
  wire[3:0] nextGrantUInt;
  wire[3:0] T139;
  wire[2:0] T140;
  wire[1:0] T141;
  wire T142;
  wire[1:0] T143;
  wire[1:0] T144;
  wire[3:0] T145;
  wire[3:0] T146;
  wire[7:0] T147;
  wire[7:0] T148;
  wire[1:0] T149;
  wire[3:0] T150;
  wire[1:0] T151;
  wire T152;
  wire T153;
  wire T154;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire[3:0] T68;
  wire[3:0] T69;
  wire T70;
  wire T71;
  wire T72;
  wire T73;
  wire[3:0] T74;
  wire[3:0] T75;
  wire T76;
  wire[1:0] T155;
  wire[3:0] T156;
  wire[1:0] T157;
  wire T158;
  wire T159;
  wire T160;
  wire T77;
  wire T78;
  wire T79;
  wire T80;
  wire T81;
  wire T82;
  wire[3:0] T83;
  wire T84;
  wire T85;
  wire T86;
  wire T87;
  wire T88;
  wire T89;
  wire T90;
  wire T91;
  wire T92;
  wire T93;
  wire T94;
  wire T95;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  wire T101;
  wire T102;
  wire T103;
  wire T104;
  wire T105;
  wire T106;
  wire T107;
  wire T108;
  wire T109;
  wire T110;
  wire T111;
  wire T112;
  wire T113;
  wire T114;
  wire T115;
  wire T116;
  wire T117;
  wire T118;
  wire T119;
  wire T120;
  wire T121;
  wire T122;
  wire T123;
  wire T124;
  wire T125;
  wire T126;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    nextGrant = {1{1'b0}};
  end
// synthesis translate_on
`endif

  assign io_chosen = T127;
  assign T127 = {T160, T128};
  assign T128 = {T159, T129};
  assign T129 = {T158, T130};
  assign T130 = T131[1'h1:1'h1];
  assign T131 = T157 | T132;
  assign T132 = T133[1'h1:1'h0];
  assign T133 = T156 | T134;
  assign T134 = T135[2'h3:1'h0];
  assign T135 = T155 | T136;
  assign T136 = winner[3'h7:1'h0];
  assign winner = T1;
  assign T1 = T41 ? T5 : nextGrant;
  assign T137 = reset ? 10'h200 : T2;
  assign T2 = T41 ? T3 : nextGrant;
  assign T3 = T4 ? winner : nextGrant;
  assign T4 = winner != 10'h0;
  assign T5 = T24 & requestsBits;
  assign requestsBits = {T15, T6};
  assign T6 = {T12, T7};
  assign T7 = {T11, T8};
  assign T8 = {T10, T9};
  assign T9 = io_requests_0_request;
  assign T10 = io_requests_1_request;
  assign T11 = io_requests_2_request;
  assign T12 = {T14, T13};
  assign T13 = io_requests_3_request;
  assign T14 = io_requests_4_request;
  assign T15 = {T21, T16};
  assign T16 = {T20, T17};
  assign T17 = {T19, T18};
  assign T18 = io_requests_5_request;
  assign T19 = io_requests_6_request;
  assign T20 = io_requests_7_request;
  assign T21 = {T23, T22};
  assign T22 = io_requests_8_request;
  assign T23 = io_requests_9_request;
  assign T24 = T40 ? passSelectL1 : T25;
  assign T25 = passSelectL0[4'h9:1'h0];
  assign passSelectL0 = T26;
  assign T26 = T41 ? T27 : 11'h0;
  assign T27 = T33 + T28;
  assign T28 = {T32, T29};
  assign T29 = {T31, T30};
  assign T30 = nextGrant[4'h9:4'h9];
  assign T31 = nextGrant[4'h8:1'h0];
  assign T32 = 1'h0;
  assign T33 = {T35, T34};
  assign T34 = ~ requestsBits;
  assign T35 = 1'h0;
  assign passSelectL1 = T36;
  assign T36 = T41 ? T37 : 10'h0;
  assign T37 = T39 + T138;
  assign T138 = {9'h0, T38};
  assign T38 = 1'h1;
  assign T39 = ~ requestsBits;
  assign T40 = passSelectL0[4'ha:4'ha];
  assign T41 = T42 ^ 1'h1;
  assign T42 = T64 & T43;
  assign T43 = ~ lockRelease;
  assign lockRelease = T44;
  assign T44 = T63 ? T61 : T45;
  assign T45 = T60 ? T54 : T46;
  assign T46 = T53 ? T51 : T47;
  assign T47 = T48 ? io_requests_1_releaseLock : io_requests_0_releaseLock;
  assign T48 = T49[1'h0:1'h0];
  assign T49 = nextGrantUInt;
  assign nextGrantUInt = T139;
  assign T139 = {T154, T140};
  assign T140 = {T153, T141};
  assign T141 = {T152, T142};
  assign T142 = T143[1'h1:1'h1];
  assign T143 = T151 | T144;
  assign T144 = T145[1'h1:1'h0];
  assign T145 = T150 | T146;
  assign T146 = T147[2'h3:1'h0];
  assign T147 = T149 | T148;
  assign T148 = nextGrant[3'h7:1'h0];
  assign T149 = nextGrant[4'h9:4'h8];
  assign T150 = T147[3'h7:3'h4];
  assign T151 = T145[2'h3:2'h2];
  assign T152 = T151 != 2'h0;
  assign T153 = T150 != 4'h0;
  assign T154 = T149 != 2'h0;
  assign T51 = T52 ? io_requests_3_releaseLock : io_requests_2_releaseLock;
  assign T52 = T49[1'h0:1'h0];
  assign T53 = T49[1'h1:1'h1];
  assign T54 = T59 ? T57 : T55;
  assign T55 = T56 ? io_requests_5_releaseLock : io_requests_4_releaseLock;
  assign T56 = T49[1'h0:1'h0];
  assign T57 = T58 ? io_requests_7_releaseLock : io_requests_6_releaseLock;
  assign T58 = T49[1'h0:1'h0];
  assign T59 = T49[1'h1:1'h1];
  assign T60 = T49[2'h2:2'h2];
  assign T61 = T62 ? io_requests_9_releaseLock : io_requests_8_releaseLock;
  assign T62 = T49[1'h0:1'h0];
  assign T63 = T49[2'h3:2'h3];
  assign T64 = T71 & T65;
  assign T65 = T70 & T66;
  assign T66 = T67 - 1'h1;
  assign T67 = 1'h1 << T68;
  assign T68 = T69 + 4'h1;
  assign T69 = nextGrantUInt - nextGrantUInt;
  assign T70 = requestsBits >> nextGrantUInt;
  assign T71 = T76 & T72;
  assign T72 = T73 - 1'h1;
  assign T73 = 1'h1 << T74;
  assign T74 = T75 + 4'h1;
  assign T75 = nextGrantUInt - nextGrantUInt;
  assign T76 = nextGrant >> nextGrantUInt;
  assign T155 = winner[4'h9:4'h8];
  assign T156 = T135[3'h7:3'h4];
  assign T157 = T133[2'h3:2'h2];
  assign T158 = T157 != 2'h0;
  assign T159 = T156 != 4'h0;
  assign T160 = T155 != 2'h0;
  assign io_resource_valid = T77;
  assign T77 = T78 & io_resource_ready;
  assign T78 = T96 ? T94 : T79;
  assign T79 = T93 ? T87 : T80;
  assign T80 = T86 ? T84 : T81;
  assign T81 = T82 ? io_requests_1_grant : io_requests_0_grant;
  assign T82 = T83[1'h0:1'h0];
  assign T83 = io_chosen;
  assign T84 = T85 ? io_requests_3_grant : io_requests_2_grant;
  assign T85 = T83[1'h0:1'h0];
  assign T86 = T83[1'h1:1'h1];
  assign T87 = T92 ? T90 : T88;
  assign T88 = T89 ? io_requests_5_grant : io_requests_4_grant;
  assign T89 = T83[1'h0:1'h0];
  assign T90 = T91 ? io_requests_7_grant : io_requests_6_grant;
  assign T91 = T83[1'h0:1'h0];
  assign T92 = T83[1'h1:1'h1];
  assign T93 = T83[2'h2:2'h2];
  assign T94 = T95 ? io_requests_9_grant : io_requests_8_grant;
  assign T95 = T83[1'h0:1'h0];
  assign T96 = T83[2'h3:2'h3];
  assign io_requests_0_grant = T97;
  assign T97 = T98 & io_resource_ready;
  assign T98 = T99;
  assign T99 = winner[1'h0:1'h0];
  assign io_requests_1_grant = T100;
  assign T100 = T101 & io_resource_ready;
  assign T101 = T102;
  assign T102 = winner[1'h1:1'h1];
  assign io_requests_2_grant = T103;
  assign T103 = T104 & io_resource_ready;
  assign T104 = T105;
  assign T105 = winner[2'h2:2'h2];
  assign io_requests_3_grant = T106;
  assign T106 = T107 & io_resource_ready;
  assign T107 = T108;
  assign T108 = winner[2'h3:2'h3];
  assign io_requests_4_grant = T109;
  assign T109 = T110 & io_resource_ready;
  assign T110 = T111;
  assign T111 = winner[3'h4:3'h4];
  assign io_requests_5_grant = T112;
  assign T112 = T113 & io_resource_ready;
  assign T113 = T114;
  assign T114 = winner[3'h5:3'h5];
  assign io_requests_6_grant = T115;
  assign T115 = T116 & io_resource_ready;
  assign T116 = T117;
  assign T117 = winner[3'h6:3'h6];
  assign io_requests_7_grant = T118;
  assign T118 = T119 & io_resource_ready;
  assign T119 = T120;
  assign T120 = winner[3'h7:3'h7];
  assign io_requests_8_grant = T121;
  assign T121 = T122 & io_resource_ready;
  assign T122 = T123;
  assign T123 = winner[4'h8:4'h8];
  assign io_requests_9_grant = T124;
  assign T124 = T125 & io_resource_ready;
  assign T125 = T126;
  assign T126 = winner[4'h9:4'h9];

  always @(posedge clk) begin
    if(reset) begin
      nextGrant <= 10'h200;
    end else if(T41) begin
      nextGrant <= T3;
    end
  end
endmodule

module SwitchAllocator_1(input clk, input reset,
    input  io_requests_9_9_releaseLock,
    output io_requests_9_9_grant,
    input  io_requests_9_9_request,
    input [2:0] io_requests_9_9_priorityLevel,
    input  io_requests_9_8_releaseLock,
    output io_requests_9_8_grant,
    input  io_requests_9_8_request,
    input [2:0] io_requests_9_8_priorityLevel,
    input  io_requests_9_7_releaseLock,
    output io_requests_9_7_grant,
    input  io_requests_9_7_request,
    input [2:0] io_requests_9_7_priorityLevel,
    input  io_requests_9_6_releaseLock,
    output io_requests_9_6_grant,
    input  io_requests_9_6_request,
    input [2:0] io_requests_9_6_priorityLevel,
    input  io_requests_9_5_releaseLock,
    output io_requests_9_5_grant,
    input  io_requests_9_5_request,
    input [2:0] io_requests_9_5_priorityLevel,
    input  io_requests_9_4_releaseLock,
    output io_requests_9_4_grant,
    input  io_requests_9_4_request,
    input [2:0] io_requests_9_4_priorityLevel,
    input  io_requests_9_3_releaseLock,
    output io_requests_9_3_grant,
    input  io_requests_9_3_request,
    input [2:0] io_requests_9_3_priorityLevel,
    input  io_requests_9_2_releaseLock,
    output io_requests_9_2_grant,
    input  io_requests_9_2_request,
    input [2:0] io_requests_9_2_priorityLevel,
    input  io_requests_9_1_releaseLock,
    output io_requests_9_1_grant,
    input  io_requests_9_1_request,
    input [2:0] io_requests_9_1_priorityLevel,
    input  io_requests_9_0_releaseLock,
    output io_requests_9_0_grant,
    input  io_requests_9_0_request,
    input [2:0] io_requests_9_0_priorityLevel,
    input  io_requests_8_9_releaseLock,
    output io_requests_8_9_grant,
    input  io_requests_8_9_request,
    input [2:0] io_requests_8_9_priorityLevel,
    input  io_requests_8_8_releaseLock,
    output io_requests_8_8_grant,
    input  io_requests_8_8_request,
    input [2:0] io_requests_8_8_priorityLevel,
    input  io_requests_8_7_releaseLock,
    output io_requests_8_7_grant,
    input  io_requests_8_7_request,
    input [2:0] io_requests_8_7_priorityLevel,
    input  io_requests_8_6_releaseLock,
    output io_requests_8_6_grant,
    input  io_requests_8_6_request,
    input [2:0] io_requests_8_6_priorityLevel,
    input  io_requests_8_5_releaseLock,
    output io_requests_8_5_grant,
    input  io_requests_8_5_request,
    input [2:0] io_requests_8_5_priorityLevel,
    input  io_requests_8_4_releaseLock,
    output io_requests_8_4_grant,
    input  io_requests_8_4_request,
    input [2:0] io_requests_8_4_priorityLevel,
    input  io_requests_8_3_releaseLock,
    output io_requests_8_3_grant,
    input  io_requests_8_3_request,
    input [2:0] io_requests_8_3_priorityLevel,
    input  io_requests_8_2_releaseLock,
    output io_requests_8_2_grant,
    input  io_requests_8_2_request,
    input [2:0] io_requests_8_2_priorityLevel,
    input  io_requests_8_1_releaseLock,
    output io_requests_8_1_grant,
    input  io_requests_8_1_request,
    input [2:0] io_requests_8_1_priorityLevel,
    input  io_requests_8_0_releaseLock,
    output io_requests_8_0_grant,
    input  io_requests_8_0_request,
    input [2:0] io_requests_8_0_priorityLevel,
    input  io_requests_7_9_releaseLock,
    output io_requests_7_9_grant,
    input  io_requests_7_9_request,
    input [2:0] io_requests_7_9_priorityLevel,
    input  io_requests_7_8_releaseLock,
    output io_requests_7_8_grant,
    input  io_requests_7_8_request,
    input [2:0] io_requests_7_8_priorityLevel,
    input  io_requests_7_7_releaseLock,
    output io_requests_7_7_grant,
    input  io_requests_7_7_request,
    input [2:0] io_requests_7_7_priorityLevel,
    input  io_requests_7_6_releaseLock,
    output io_requests_7_6_grant,
    input  io_requests_7_6_request,
    input [2:0] io_requests_7_6_priorityLevel,
    input  io_requests_7_5_releaseLock,
    output io_requests_7_5_grant,
    input  io_requests_7_5_request,
    input [2:0] io_requests_7_5_priorityLevel,
    input  io_requests_7_4_releaseLock,
    output io_requests_7_4_grant,
    input  io_requests_7_4_request,
    input [2:0] io_requests_7_4_priorityLevel,
    input  io_requests_7_3_releaseLock,
    output io_requests_7_3_grant,
    input  io_requests_7_3_request,
    input [2:0] io_requests_7_3_priorityLevel,
    input  io_requests_7_2_releaseLock,
    output io_requests_7_2_grant,
    input  io_requests_7_2_request,
    input [2:0] io_requests_7_2_priorityLevel,
    input  io_requests_7_1_releaseLock,
    output io_requests_7_1_grant,
    input  io_requests_7_1_request,
    input [2:0] io_requests_7_1_priorityLevel,
    input  io_requests_7_0_releaseLock,
    output io_requests_7_0_grant,
    input  io_requests_7_0_request,
    input [2:0] io_requests_7_0_priorityLevel,
    input  io_requests_6_9_releaseLock,
    output io_requests_6_9_grant,
    input  io_requests_6_9_request,
    input [2:0] io_requests_6_9_priorityLevel,
    input  io_requests_6_8_releaseLock,
    output io_requests_6_8_grant,
    input  io_requests_6_8_request,
    input [2:0] io_requests_6_8_priorityLevel,
    input  io_requests_6_7_releaseLock,
    output io_requests_6_7_grant,
    input  io_requests_6_7_request,
    input [2:0] io_requests_6_7_priorityLevel,
    input  io_requests_6_6_releaseLock,
    output io_requests_6_6_grant,
    input  io_requests_6_6_request,
    input [2:0] io_requests_6_6_priorityLevel,
    input  io_requests_6_5_releaseLock,
    output io_requests_6_5_grant,
    input  io_requests_6_5_request,
    input [2:0] io_requests_6_5_priorityLevel,
    input  io_requests_6_4_releaseLock,
    output io_requests_6_4_grant,
    input  io_requests_6_4_request,
    input [2:0] io_requests_6_4_priorityLevel,
    input  io_requests_6_3_releaseLock,
    output io_requests_6_3_grant,
    input  io_requests_6_3_request,
    input [2:0] io_requests_6_3_priorityLevel,
    input  io_requests_6_2_releaseLock,
    output io_requests_6_2_grant,
    input  io_requests_6_2_request,
    input [2:0] io_requests_6_2_priorityLevel,
    input  io_requests_6_1_releaseLock,
    output io_requests_6_1_grant,
    input  io_requests_6_1_request,
    input [2:0] io_requests_6_1_priorityLevel,
    input  io_requests_6_0_releaseLock,
    output io_requests_6_0_grant,
    input  io_requests_6_0_request,
    input [2:0] io_requests_6_0_priorityLevel,
    input  io_requests_5_9_releaseLock,
    output io_requests_5_9_grant,
    input  io_requests_5_9_request,
    input [2:0] io_requests_5_9_priorityLevel,
    input  io_requests_5_8_releaseLock,
    output io_requests_5_8_grant,
    input  io_requests_5_8_request,
    input [2:0] io_requests_5_8_priorityLevel,
    input  io_requests_5_7_releaseLock,
    output io_requests_5_7_grant,
    input  io_requests_5_7_request,
    input [2:0] io_requests_5_7_priorityLevel,
    input  io_requests_5_6_releaseLock,
    output io_requests_5_6_grant,
    input  io_requests_5_6_request,
    input [2:0] io_requests_5_6_priorityLevel,
    input  io_requests_5_5_releaseLock,
    output io_requests_5_5_grant,
    input  io_requests_5_5_request,
    input [2:0] io_requests_5_5_priorityLevel,
    input  io_requests_5_4_releaseLock,
    output io_requests_5_4_grant,
    input  io_requests_5_4_request,
    input [2:0] io_requests_5_4_priorityLevel,
    input  io_requests_5_3_releaseLock,
    output io_requests_5_3_grant,
    input  io_requests_5_3_request,
    input [2:0] io_requests_5_3_priorityLevel,
    input  io_requests_5_2_releaseLock,
    output io_requests_5_2_grant,
    input  io_requests_5_2_request,
    input [2:0] io_requests_5_2_priorityLevel,
    input  io_requests_5_1_releaseLock,
    output io_requests_5_1_grant,
    input  io_requests_5_1_request,
    input [2:0] io_requests_5_1_priorityLevel,
    input  io_requests_5_0_releaseLock,
    output io_requests_5_0_grant,
    input  io_requests_5_0_request,
    input [2:0] io_requests_5_0_priorityLevel,
    input  io_requests_4_9_releaseLock,
    output io_requests_4_9_grant,
    input  io_requests_4_9_request,
    input [2:0] io_requests_4_9_priorityLevel,
    input  io_requests_4_8_releaseLock,
    output io_requests_4_8_grant,
    input  io_requests_4_8_request,
    input [2:0] io_requests_4_8_priorityLevel,
    input  io_requests_4_7_releaseLock,
    output io_requests_4_7_grant,
    input  io_requests_4_7_request,
    input [2:0] io_requests_4_7_priorityLevel,
    input  io_requests_4_6_releaseLock,
    output io_requests_4_6_grant,
    input  io_requests_4_6_request,
    input [2:0] io_requests_4_6_priorityLevel,
    input  io_requests_4_5_releaseLock,
    output io_requests_4_5_grant,
    input  io_requests_4_5_request,
    input [2:0] io_requests_4_5_priorityLevel,
    input  io_requests_4_4_releaseLock,
    output io_requests_4_4_grant,
    input  io_requests_4_4_request,
    input [2:0] io_requests_4_4_priorityLevel,
    input  io_requests_4_3_releaseLock,
    output io_requests_4_3_grant,
    input  io_requests_4_3_request,
    input [2:0] io_requests_4_3_priorityLevel,
    input  io_requests_4_2_releaseLock,
    output io_requests_4_2_grant,
    input  io_requests_4_2_request,
    input [2:0] io_requests_4_2_priorityLevel,
    input  io_requests_4_1_releaseLock,
    output io_requests_4_1_grant,
    input  io_requests_4_1_request,
    input [2:0] io_requests_4_1_priorityLevel,
    input  io_requests_4_0_releaseLock,
    output io_requests_4_0_grant,
    input  io_requests_4_0_request,
    input [2:0] io_requests_4_0_priorityLevel,
    input  io_requests_3_9_releaseLock,
    output io_requests_3_9_grant,
    input  io_requests_3_9_request,
    input [2:0] io_requests_3_9_priorityLevel,
    input  io_requests_3_8_releaseLock,
    output io_requests_3_8_grant,
    input  io_requests_3_8_request,
    input [2:0] io_requests_3_8_priorityLevel,
    input  io_requests_3_7_releaseLock,
    output io_requests_3_7_grant,
    input  io_requests_3_7_request,
    input [2:0] io_requests_3_7_priorityLevel,
    input  io_requests_3_6_releaseLock,
    output io_requests_3_6_grant,
    input  io_requests_3_6_request,
    input [2:0] io_requests_3_6_priorityLevel,
    input  io_requests_3_5_releaseLock,
    output io_requests_3_5_grant,
    input  io_requests_3_5_request,
    input [2:0] io_requests_3_5_priorityLevel,
    input  io_requests_3_4_releaseLock,
    output io_requests_3_4_grant,
    input  io_requests_3_4_request,
    input [2:0] io_requests_3_4_priorityLevel,
    input  io_requests_3_3_releaseLock,
    output io_requests_3_3_grant,
    input  io_requests_3_3_request,
    input [2:0] io_requests_3_3_priorityLevel,
    input  io_requests_3_2_releaseLock,
    output io_requests_3_2_grant,
    input  io_requests_3_2_request,
    input [2:0] io_requests_3_2_priorityLevel,
    input  io_requests_3_1_releaseLock,
    output io_requests_3_1_grant,
    input  io_requests_3_1_request,
    input [2:0] io_requests_3_1_priorityLevel,
    input  io_requests_3_0_releaseLock,
    output io_requests_3_0_grant,
    input  io_requests_3_0_request,
    input [2:0] io_requests_3_0_priorityLevel,
    input  io_requests_2_9_releaseLock,
    output io_requests_2_9_grant,
    input  io_requests_2_9_request,
    input [2:0] io_requests_2_9_priorityLevel,
    input  io_requests_2_8_releaseLock,
    output io_requests_2_8_grant,
    input  io_requests_2_8_request,
    input [2:0] io_requests_2_8_priorityLevel,
    input  io_requests_2_7_releaseLock,
    output io_requests_2_7_grant,
    input  io_requests_2_7_request,
    input [2:0] io_requests_2_7_priorityLevel,
    input  io_requests_2_6_releaseLock,
    output io_requests_2_6_grant,
    input  io_requests_2_6_request,
    input [2:0] io_requests_2_6_priorityLevel,
    input  io_requests_2_5_releaseLock,
    output io_requests_2_5_grant,
    input  io_requests_2_5_request,
    input [2:0] io_requests_2_5_priorityLevel,
    input  io_requests_2_4_releaseLock,
    output io_requests_2_4_grant,
    input  io_requests_2_4_request,
    input [2:0] io_requests_2_4_priorityLevel,
    input  io_requests_2_3_releaseLock,
    output io_requests_2_3_grant,
    input  io_requests_2_3_request,
    input [2:0] io_requests_2_3_priorityLevel,
    input  io_requests_2_2_releaseLock,
    output io_requests_2_2_grant,
    input  io_requests_2_2_request,
    input [2:0] io_requests_2_2_priorityLevel,
    input  io_requests_2_1_releaseLock,
    output io_requests_2_1_grant,
    input  io_requests_2_1_request,
    input [2:0] io_requests_2_1_priorityLevel,
    input  io_requests_2_0_releaseLock,
    output io_requests_2_0_grant,
    input  io_requests_2_0_request,
    input [2:0] io_requests_2_0_priorityLevel,
    input  io_requests_1_9_releaseLock,
    output io_requests_1_9_grant,
    input  io_requests_1_9_request,
    input [2:0] io_requests_1_9_priorityLevel,
    input  io_requests_1_8_releaseLock,
    output io_requests_1_8_grant,
    input  io_requests_1_8_request,
    input [2:0] io_requests_1_8_priorityLevel,
    input  io_requests_1_7_releaseLock,
    output io_requests_1_7_grant,
    input  io_requests_1_7_request,
    input [2:0] io_requests_1_7_priorityLevel,
    input  io_requests_1_6_releaseLock,
    output io_requests_1_6_grant,
    input  io_requests_1_6_request,
    input [2:0] io_requests_1_6_priorityLevel,
    input  io_requests_1_5_releaseLock,
    output io_requests_1_5_grant,
    input  io_requests_1_5_request,
    input [2:0] io_requests_1_5_priorityLevel,
    input  io_requests_1_4_releaseLock,
    output io_requests_1_4_grant,
    input  io_requests_1_4_request,
    input [2:0] io_requests_1_4_priorityLevel,
    input  io_requests_1_3_releaseLock,
    output io_requests_1_3_grant,
    input  io_requests_1_3_request,
    input [2:0] io_requests_1_3_priorityLevel,
    input  io_requests_1_2_releaseLock,
    output io_requests_1_2_grant,
    input  io_requests_1_2_request,
    input [2:0] io_requests_1_2_priorityLevel,
    input  io_requests_1_1_releaseLock,
    output io_requests_1_1_grant,
    input  io_requests_1_1_request,
    input [2:0] io_requests_1_1_priorityLevel,
    input  io_requests_1_0_releaseLock,
    output io_requests_1_0_grant,
    input  io_requests_1_0_request,
    input [2:0] io_requests_1_0_priorityLevel,
    input  io_requests_0_9_releaseLock,
    output io_requests_0_9_grant,
    input  io_requests_0_9_request,
    input [2:0] io_requests_0_9_priorityLevel,
    input  io_requests_0_8_releaseLock,
    output io_requests_0_8_grant,
    input  io_requests_0_8_request,
    input [2:0] io_requests_0_8_priorityLevel,
    input  io_requests_0_7_releaseLock,
    output io_requests_0_7_grant,
    input  io_requests_0_7_request,
    input [2:0] io_requests_0_7_priorityLevel,
    input  io_requests_0_6_releaseLock,
    output io_requests_0_6_grant,
    input  io_requests_0_6_request,
    input [2:0] io_requests_0_6_priorityLevel,
    input  io_requests_0_5_releaseLock,
    output io_requests_0_5_grant,
    input  io_requests_0_5_request,
    input [2:0] io_requests_0_5_priorityLevel,
    input  io_requests_0_4_releaseLock,
    output io_requests_0_4_grant,
    input  io_requests_0_4_request,
    input [2:0] io_requests_0_4_priorityLevel,
    input  io_requests_0_3_releaseLock,
    output io_requests_0_3_grant,
    input  io_requests_0_3_request,
    input [2:0] io_requests_0_3_priorityLevel,
    input  io_requests_0_2_releaseLock,
    output io_requests_0_2_grant,
    input  io_requests_0_2_request,
    input [2:0] io_requests_0_2_priorityLevel,
    input  io_requests_0_1_releaseLock,
    output io_requests_0_1_grant,
    input  io_requests_0_1_request,
    input [2:0] io_requests_0_1_priorityLevel,
    input  io_requests_0_0_releaseLock,
    output io_requests_0_0_grant,
    input  io_requests_0_0_request,
    input [2:0] io_requests_0_0_priorityLevel,
    input  io_resources_9_ready,
    output io_resources_9_valid,
    input  io_resources_8_ready,
    output io_resources_8_valid,
    input  io_resources_7_ready,
    output io_resources_7_valid,
    input  io_resources_6_ready,
    output io_resources_6_valid,
    input  io_resources_5_ready,
    output io_resources_5_valid,
    input  io_resources_4_ready,
    output io_resources_4_valid,
    input  io_resources_3_ready,
    output io_resources_3_valid,
    input  io_resources_2_ready,
    output io_resources_2_valid,
    input  io_resources_1_ready,
    output io_resources_1_valid,
    input  io_resources_0_ready,
    output io_resources_0_valid,
    output[3:0] io_chosens_9,
    output[3:0] io_chosens_8,
    output[3:0] io_chosens_7,
    output[3:0] io_chosens_6,
    output[3:0] io_chosens_5,
    output[3:0] io_chosens_4,
    output[3:0] io_chosens_3,
    output[3:0] io_chosens_2,
    output[3:0] io_chosens_1,
    output[3:0] io_chosens_0
);

  wire RRArbiter_io_requests_9_grant;
  wire RRArbiter_io_requests_8_grant;
  wire RRArbiter_io_requests_7_grant;
  wire RRArbiter_io_requests_6_grant;
  wire RRArbiter_io_requests_5_grant;
  wire RRArbiter_io_requests_4_grant;
  wire RRArbiter_io_requests_3_grant;
  wire RRArbiter_io_requests_2_grant;
  wire RRArbiter_io_requests_1_grant;
  wire RRArbiter_io_requests_0_grant;
  wire RRArbiter_io_resource_valid;
  wire[3:0] RRArbiter_io_chosen;
  wire RRArbiter_1_io_requests_9_grant;
  wire RRArbiter_1_io_requests_8_grant;
  wire RRArbiter_1_io_requests_7_grant;
  wire RRArbiter_1_io_requests_6_grant;
  wire RRArbiter_1_io_requests_5_grant;
  wire RRArbiter_1_io_requests_4_grant;
  wire RRArbiter_1_io_requests_3_grant;
  wire RRArbiter_1_io_requests_2_grant;
  wire RRArbiter_1_io_requests_1_grant;
  wire RRArbiter_1_io_requests_0_grant;
  wire RRArbiter_1_io_resource_valid;
  wire[3:0] RRArbiter_1_io_chosen;
  wire RRArbiter_2_io_requests_9_grant;
  wire RRArbiter_2_io_requests_8_grant;
  wire RRArbiter_2_io_requests_7_grant;
  wire RRArbiter_2_io_requests_6_grant;
  wire RRArbiter_2_io_requests_5_grant;
  wire RRArbiter_2_io_requests_4_grant;
  wire RRArbiter_2_io_requests_3_grant;
  wire RRArbiter_2_io_requests_2_grant;
  wire RRArbiter_2_io_requests_1_grant;
  wire RRArbiter_2_io_requests_0_grant;
  wire RRArbiter_2_io_resource_valid;
  wire[3:0] RRArbiter_2_io_chosen;
  wire RRArbiter_3_io_requests_9_grant;
  wire RRArbiter_3_io_requests_8_grant;
  wire RRArbiter_3_io_requests_7_grant;
  wire RRArbiter_3_io_requests_6_grant;
  wire RRArbiter_3_io_requests_5_grant;
  wire RRArbiter_3_io_requests_4_grant;
  wire RRArbiter_3_io_requests_3_grant;
  wire RRArbiter_3_io_requests_2_grant;
  wire RRArbiter_3_io_requests_1_grant;
  wire RRArbiter_3_io_requests_0_grant;
  wire RRArbiter_3_io_resource_valid;
  wire[3:0] RRArbiter_3_io_chosen;
  wire RRArbiter_4_io_requests_9_grant;
  wire RRArbiter_4_io_requests_8_grant;
  wire RRArbiter_4_io_requests_7_grant;
  wire RRArbiter_4_io_requests_6_grant;
  wire RRArbiter_4_io_requests_5_grant;
  wire RRArbiter_4_io_requests_4_grant;
  wire RRArbiter_4_io_requests_3_grant;
  wire RRArbiter_4_io_requests_2_grant;
  wire RRArbiter_4_io_requests_1_grant;
  wire RRArbiter_4_io_requests_0_grant;
  wire RRArbiter_4_io_resource_valid;
  wire[3:0] RRArbiter_4_io_chosen;
  wire RRArbiter_5_io_requests_9_grant;
  wire RRArbiter_5_io_requests_8_grant;
  wire RRArbiter_5_io_requests_7_grant;
  wire RRArbiter_5_io_requests_6_grant;
  wire RRArbiter_5_io_requests_5_grant;
  wire RRArbiter_5_io_requests_4_grant;
  wire RRArbiter_5_io_requests_3_grant;
  wire RRArbiter_5_io_requests_2_grant;
  wire RRArbiter_5_io_requests_1_grant;
  wire RRArbiter_5_io_requests_0_grant;
  wire RRArbiter_5_io_resource_valid;
  wire[3:0] RRArbiter_5_io_chosen;
  wire RRArbiter_6_io_requests_9_grant;
  wire RRArbiter_6_io_requests_8_grant;
  wire RRArbiter_6_io_requests_7_grant;
  wire RRArbiter_6_io_requests_6_grant;
  wire RRArbiter_6_io_requests_5_grant;
  wire RRArbiter_6_io_requests_4_grant;
  wire RRArbiter_6_io_requests_3_grant;
  wire RRArbiter_6_io_requests_2_grant;
  wire RRArbiter_6_io_requests_1_grant;
  wire RRArbiter_6_io_requests_0_grant;
  wire RRArbiter_6_io_resource_valid;
  wire[3:0] RRArbiter_6_io_chosen;
  wire RRArbiter_7_io_requests_9_grant;
  wire RRArbiter_7_io_requests_8_grant;
  wire RRArbiter_7_io_requests_7_grant;
  wire RRArbiter_7_io_requests_6_grant;
  wire RRArbiter_7_io_requests_5_grant;
  wire RRArbiter_7_io_requests_4_grant;
  wire RRArbiter_7_io_requests_3_grant;
  wire RRArbiter_7_io_requests_2_grant;
  wire RRArbiter_7_io_requests_1_grant;
  wire RRArbiter_7_io_requests_0_grant;
  wire RRArbiter_7_io_resource_valid;
  wire[3:0] RRArbiter_7_io_chosen;
  wire RRArbiter_8_io_requests_9_grant;
  wire RRArbiter_8_io_requests_8_grant;
  wire RRArbiter_8_io_requests_7_grant;
  wire RRArbiter_8_io_requests_6_grant;
  wire RRArbiter_8_io_requests_5_grant;
  wire RRArbiter_8_io_requests_4_grant;
  wire RRArbiter_8_io_requests_3_grant;
  wire RRArbiter_8_io_requests_2_grant;
  wire RRArbiter_8_io_requests_1_grant;
  wire RRArbiter_8_io_requests_0_grant;
  wire RRArbiter_8_io_resource_valid;
  wire[3:0] RRArbiter_8_io_chosen;
  wire RRArbiter_9_io_requests_9_grant;
  wire RRArbiter_9_io_requests_8_grant;
  wire RRArbiter_9_io_requests_7_grant;
  wire RRArbiter_9_io_requests_6_grant;
  wire RRArbiter_9_io_requests_5_grant;
  wire RRArbiter_9_io_requests_4_grant;
  wire RRArbiter_9_io_requests_3_grant;
  wire RRArbiter_9_io_requests_2_grant;
  wire RRArbiter_9_io_requests_1_grant;
  wire RRArbiter_9_io_requests_0_grant;
  wire RRArbiter_9_io_resource_valid;
  wire[3:0] RRArbiter_9_io_chosen;


  assign io_chosens_0 = RRArbiter_io_chosen;
  assign io_chosens_1 = RRArbiter_1_io_chosen;
  assign io_chosens_2 = RRArbiter_2_io_chosen;
  assign io_chosens_3 = RRArbiter_3_io_chosen;
  assign io_chosens_4 = RRArbiter_4_io_chosen;
  assign io_chosens_5 = RRArbiter_5_io_chosen;
  assign io_chosens_6 = RRArbiter_6_io_chosen;
  assign io_chosens_7 = RRArbiter_7_io_chosen;
  assign io_chosens_8 = RRArbiter_8_io_chosen;
  assign io_chosens_9 = RRArbiter_9_io_chosen;
  assign io_resources_0_valid = RRArbiter_io_resource_valid;
  assign io_resources_1_valid = RRArbiter_1_io_resource_valid;
  assign io_resources_2_valid = RRArbiter_2_io_resource_valid;
  assign io_resources_3_valid = RRArbiter_3_io_resource_valid;
  assign io_resources_4_valid = RRArbiter_4_io_resource_valid;
  assign io_resources_5_valid = RRArbiter_5_io_resource_valid;
  assign io_resources_6_valid = RRArbiter_6_io_resource_valid;
  assign io_resources_7_valid = RRArbiter_7_io_resource_valid;
  assign io_resources_8_valid = RRArbiter_8_io_resource_valid;
  assign io_resources_9_valid = RRArbiter_9_io_resource_valid;
  assign io_requests_0_0_grant = RRArbiter_io_requests_0_grant;
  assign io_requests_0_1_grant = RRArbiter_io_requests_1_grant;
  assign io_requests_0_2_grant = RRArbiter_io_requests_2_grant;
  assign io_requests_0_3_grant = RRArbiter_io_requests_3_grant;
  assign io_requests_0_4_grant = RRArbiter_io_requests_4_grant;
  assign io_requests_0_5_grant = RRArbiter_io_requests_5_grant;
  assign io_requests_0_6_grant = RRArbiter_io_requests_6_grant;
  assign io_requests_0_7_grant = RRArbiter_io_requests_7_grant;
  assign io_requests_0_8_grant = RRArbiter_io_requests_8_grant;
  assign io_requests_0_9_grant = RRArbiter_io_requests_9_grant;
  assign io_requests_1_0_grant = RRArbiter_1_io_requests_0_grant;
  assign io_requests_1_1_grant = RRArbiter_1_io_requests_1_grant;
  assign io_requests_1_2_grant = RRArbiter_1_io_requests_2_grant;
  assign io_requests_1_3_grant = RRArbiter_1_io_requests_3_grant;
  assign io_requests_1_4_grant = RRArbiter_1_io_requests_4_grant;
  assign io_requests_1_5_grant = RRArbiter_1_io_requests_5_grant;
  assign io_requests_1_6_grant = RRArbiter_1_io_requests_6_grant;
  assign io_requests_1_7_grant = RRArbiter_1_io_requests_7_grant;
  assign io_requests_1_8_grant = RRArbiter_1_io_requests_8_grant;
  assign io_requests_1_9_grant = RRArbiter_1_io_requests_9_grant;
  assign io_requests_2_0_grant = RRArbiter_2_io_requests_0_grant;
  assign io_requests_2_1_grant = RRArbiter_2_io_requests_1_grant;
  assign io_requests_2_2_grant = RRArbiter_2_io_requests_2_grant;
  assign io_requests_2_3_grant = RRArbiter_2_io_requests_3_grant;
  assign io_requests_2_4_grant = RRArbiter_2_io_requests_4_grant;
  assign io_requests_2_5_grant = RRArbiter_2_io_requests_5_grant;
  assign io_requests_2_6_grant = RRArbiter_2_io_requests_6_grant;
  assign io_requests_2_7_grant = RRArbiter_2_io_requests_7_grant;
  assign io_requests_2_8_grant = RRArbiter_2_io_requests_8_grant;
  assign io_requests_2_9_grant = RRArbiter_2_io_requests_9_grant;
  assign io_requests_3_0_grant = RRArbiter_3_io_requests_0_grant;
  assign io_requests_3_1_grant = RRArbiter_3_io_requests_1_grant;
  assign io_requests_3_2_grant = RRArbiter_3_io_requests_2_grant;
  assign io_requests_3_3_grant = RRArbiter_3_io_requests_3_grant;
  assign io_requests_3_4_grant = RRArbiter_3_io_requests_4_grant;
  assign io_requests_3_5_grant = RRArbiter_3_io_requests_5_grant;
  assign io_requests_3_6_grant = RRArbiter_3_io_requests_6_grant;
  assign io_requests_3_7_grant = RRArbiter_3_io_requests_7_grant;
  assign io_requests_3_8_grant = RRArbiter_3_io_requests_8_grant;
  assign io_requests_3_9_grant = RRArbiter_3_io_requests_9_grant;
  assign io_requests_4_0_grant = RRArbiter_4_io_requests_0_grant;
  assign io_requests_4_1_grant = RRArbiter_4_io_requests_1_grant;
  assign io_requests_4_2_grant = RRArbiter_4_io_requests_2_grant;
  assign io_requests_4_3_grant = RRArbiter_4_io_requests_3_grant;
  assign io_requests_4_4_grant = RRArbiter_4_io_requests_4_grant;
  assign io_requests_4_5_grant = RRArbiter_4_io_requests_5_grant;
  assign io_requests_4_6_grant = RRArbiter_4_io_requests_6_grant;
  assign io_requests_4_7_grant = RRArbiter_4_io_requests_7_grant;
  assign io_requests_4_8_grant = RRArbiter_4_io_requests_8_grant;
  assign io_requests_4_9_grant = RRArbiter_4_io_requests_9_grant;
  assign io_requests_5_0_grant = RRArbiter_5_io_requests_0_grant;
  assign io_requests_5_1_grant = RRArbiter_5_io_requests_1_grant;
  assign io_requests_5_2_grant = RRArbiter_5_io_requests_2_grant;
  assign io_requests_5_3_grant = RRArbiter_5_io_requests_3_grant;
  assign io_requests_5_4_grant = RRArbiter_5_io_requests_4_grant;
  assign io_requests_5_5_grant = RRArbiter_5_io_requests_5_grant;
  assign io_requests_5_6_grant = RRArbiter_5_io_requests_6_grant;
  assign io_requests_5_7_grant = RRArbiter_5_io_requests_7_grant;
  assign io_requests_5_8_grant = RRArbiter_5_io_requests_8_grant;
  assign io_requests_5_9_grant = RRArbiter_5_io_requests_9_grant;
  assign io_requests_6_0_grant = RRArbiter_6_io_requests_0_grant;
  assign io_requests_6_1_grant = RRArbiter_6_io_requests_1_grant;
  assign io_requests_6_2_grant = RRArbiter_6_io_requests_2_grant;
  assign io_requests_6_3_grant = RRArbiter_6_io_requests_3_grant;
  assign io_requests_6_4_grant = RRArbiter_6_io_requests_4_grant;
  assign io_requests_6_5_grant = RRArbiter_6_io_requests_5_grant;
  assign io_requests_6_6_grant = RRArbiter_6_io_requests_6_grant;
  assign io_requests_6_7_grant = RRArbiter_6_io_requests_7_grant;
  assign io_requests_6_8_grant = RRArbiter_6_io_requests_8_grant;
  assign io_requests_6_9_grant = RRArbiter_6_io_requests_9_grant;
  assign io_requests_7_0_grant = RRArbiter_7_io_requests_0_grant;
  assign io_requests_7_1_grant = RRArbiter_7_io_requests_1_grant;
  assign io_requests_7_2_grant = RRArbiter_7_io_requests_2_grant;
  assign io_requests_7_3_grant = RRArbiter_7_io_requests_3_grant;
  assign io_requests_7_4_grant = RRArbiter_7_io_requests_4_grant;
  assign io_requests_7_5_grant = RRArbiter_7_io_requests_5_grant;
  assign io_requests_7_6_grant = RRArbiter_7_io_requests_6_grant;
  assign io_requests_7_7_grant = RRArbiter_7_io_requests_7_grant;
  assign io_requests_7_8_grant = RRArbiter_7_io_requests_8_grant;
  assign io_requests_7_9_grant = RRArbiter_7_io_requests_9_grant;
  assign io_requests_8_0_grant = RRArbiter_8_io_requests_0_grant;
  assign io_requests_8_1_grant = RRArbiter_8_io_requests_1_grant;
  assign io_requests_8_2_grant = RRArbiter_8_io_requests_2_grant;
  assign io_requests_8_3_grant = RRArbiter_8_io_requests_3_grant;
  assign io_requests_8_4_grant = RRArbiter_8_io_requests_4_grant;
  assign io_requests_8_5_grant = RRArbiter_8_io_requests_5_grant;
  assign io_requests_8_6_grant = RRArbiter_8_io_requests_6_grant;
  assign io_requests_8_7_grant = RRArbiter_8_io_requests_7_grant;
  assign io_requests_8_8_grant = RRArbiter_8_io_requests_8_grant;
  assign io_requests_8_9_grant = RRArbiter_8_io_requests_9_grant;
  assign io_requests_9_0_grant = RRArbiter_9_io_requests_0_grant;
  assign io_requests_9_1_grant = RRArbiter_9_io_requests_1_grant;
  assign io_requests_9_2_grant = RRArbiter_9_io_requests_2_grant;
  assign io_requests_9_3_grant = RRArbiter_9_io_requests_3_grant;
  assign io_requests_9_4_grant = RRArbiter_9_io_requests_4_grant;
  assign io_requests_9_5_grant = RRArbiter_9_io_requests_5_grant;
  assign io_requests_9_6_grant = RRArbiter_9_io_requests_6_grant;
  assign io_requests_9_7_grant = RRArbiter_9_io_requests_7_grant;
  assign io_requests_9_8_grant = RRArbiter_9_io_requests_8_grant;
  assign io_requests_9_9_grant = RRArbiter_9_io_requests_9_grant;
  RRArbiter_1 RRArbiter(.clk(clk), .reset(reset),
       .io_requests_9_releaseLock( io_requests_0_9_releaseLock ),
       .io_requests_9_grant( RRArbiter_io_requests_9_grant ),
       .io_requests_9_request( io_requests_0_9_request ),
       .io_requests_9_priorityLevel( io_requests_0_9_priorityLevel ),
       .io_requests_8_releaseLock( io_requests_0_8_releaseLock ),
       .io_requests_8_grant( RRArbiter_io_requests_8_grant ),
       .io_requests_8_request( io_requests_0_8_request ),
       .io_requests_8_priorityLevel( io_requests_0_8_priorityLevel ),
       .io_requests_7_releaseLock( io_requests_0_7_releaseLock ),
       .io_requests_7_grant( RRArbiter_io_requests_7_grant ),
       .io_requests_7_request( io_requests_0_7_request ),
       .io_requests_7_priorityLevel( io_requests_0_7_priorityLevel ),
       .io_requests_6_releaseLock( io_requests_0_6_releaseLock ),
       .io_requests_6_grant( RRArbiter_io_requests_6_grant ),
       .io_requests_6_request( io_requests_0_6_request ),
       .io_requests_6_priorityLevel( io_requests_0_6_priorityLevel ),
       .io_requests_5_releaseLock( io_requests_0_5_releaseLock ),
       .io_requests_5_grant( RRArbiter_io_requests_5_grant ),
       .io_requests_5_request( io_requests_0_5_request ),
       .io_requests_5_priorityLevel( io_requests_0_5_priorityLevel ),
       .io_requests_4_releaseLock( io_requests_0_4_releaseLock ),
       .io_requests_4_grant( RRArbiter_io_requests_4_grant ),
       .io_requests_4_request( io_requests_0_4_request ),
       .io_requests_4_priorityLevel( io_requests_0_4_priorityLevel ),
       .io_requests_3_releaseLock( io_requests_0_3_releaseLock ),
       .io_requests_3_grant( RRArbiter_io_requests_3_grant ),
       .io_requests_3_request( io_requests_0_3_request ),
       .io_requests_3_priorityLevel( io_requests_0_3_priorityLevel ),
       .io_requests_2_releaseLock( io_requests_0_2_releaseLock ),
       .io_requests_2_grant( RRArbiter_io_requests_2_grant ),
       .io_requests_2_request( io_requests_0_2_request ),
       .io_requests_2_priorityLevel( io_requests_0_2_priorityLevel ),
       .io_requests_1_releaseLock( io_requests_0_1_releaseLock ),
       .io_requests_1_grant( RRArbiter_io_requests_1_grant ),
       .io_requests_1_request( io_requests_0_1_request ),
       .io_requests_1_priorityLevel( io_requests_0_1_priorityLevel ),
       .io_requests_0_releaseLock( io_requests_0_0_releaseLock ),
       .io_requests_0_grant( RRArbiter_io_requests_0_grant ),
       .io_requests_0_request( io_requests_0_0_request ),
       .io_requests_0_priorityLevel( io_requests_0_0_priorityLevel ),
       .io_resource_ready( io_resources_0_ready ),
       .io_resource_valid( RRArbiter_io_resource_valid ),
       .io_chosen( RRArbiter_io_chosen )
  );
  RRArbiter_1 RRArbiter_1(.clk(clk), .reset(reset),
       .io_requests_9_releaseLock( io_requests_1_9_releaseLock ),
       .io_requests_9_grant( RRArbiter_1_io_requests_9_grant ),
       .io_requests_9_request( io_requests_1_9_request ),
       .io_requests_9_priorityLevel( io_requests_1_9_priorityLevel ),
       .io_requests_8_releaseLock( io_requests_1_8_releaseLock ),
       .io_requests_8_grant( RRArbiter_1_io_requests_8_grant ),
       .io_requests_8_request( io_requests_1_8_request ),
       .io_requests_8_priorityLevel( io_requests_1_8_priorityLevel ),
       .io_requests_7_releaseLock( io_requests_1_7_releaseLock ),
       .io_requests_7_grant( RRArbiter_1_io_requests_7_grant ),
       .io_requests_7_request( io_requests_1_7_request ),
       .io_requests_7_priorityLevel( io_requests_1_7_priorityLevel ),
       .io_requests_6_releaseLock( io_requests_1_6_releaseLock ),
       .io_requests_6_grant( RRArbiter_1_io_requests_6_grant ),
       .io_requests_6_request( io_requests_1_6_request ),
       .io_requests_6_priorityLevel( io_requests_1_6_priorityLevel ),
       .io_requests_5_releaseLock( io_requests_1_5_releaseLock ),
       .io_requests_5_grant( RRArbiter_1_io_requests_5_grant ),
       .io_requests_5_request( io_requests_1_5_request ),
       .io_requests_5_priorityLevel( io_requests_1_5_priorityLevel ),
       .io_requests_4_releaseLock( io_requests_1_4_releaseLock ),
       .io_requests_4_grant( RRArbiter_1_io_requests_4_grant ),
       .io_requests_4_request( io_requests_1_4_request ),
       .io_requests_4_priorityLevel( io_requests_1_4_priorityLevel ),
       .io_requests_3_releaseLock( io_requests_1_3_releaseLock ),
       .io_requests_3_grant( RRArbiter_1_io_requests_3_grant ),
       .io_requests_3_request( io_requests_1_3_request ),
       .io_requests_3_priorityLevel( io_requests_1_3_priorityLevel ),
       .io_requests_2_releaseLock( io_requests_1_2_releaseLock ),
       .io_requests_2_grant( RRArbiter_1_io_requests_2_grant ),
       .io_requests_2_request( io_requests_1_2_request ),
       .io_requests_2_priorityLevel( io_requests_1_2_priorityLevel ),
       .io_requests_1_releaseLock( io_requests_1_1_releaseLock ),
       .io_requests_1_grant( RRArbiter_1_io_requests_1_grant ),
       .io_requests_1_request( io_requests_1_1_request ),
       .io_requests_1_priorityLevel( io_requests_1_1_priorityLevel ),
       .io_requests_0_releaseLock( io_requests_1_0_releaseLock ),
       .io_requests_0_grant( RRArbiter_1_io_requests_0_grant ),
       .io_requests_0_request( io_requests_1_0_request ),
       .io_requests_0_priorityLevel( io_requests_1_0_priorityLevel ),
       .io_resource_ready( io_resources_1_ready ),
       .io_resource_valid( RRArbiter_1_io_resource_valid ),
       .io_chosen( RRArbiter_1_io_chosen )
  );
  RRArbiter_1 RRArbiter_2(.clk(clk), .reset(reset),
       .io_requests_9_releaseLock( io_requests_2_9_releaseLock ),
       .io_requests_9_grant( RRArbiter_2_io_requests_9_grant ),
       .io_requests_9_request( io_requests_2_9_request ),
       .io_requests_9_priorityLevel( io_requests_2_9_priorityLevel ),
       .io_requests_8_releaseLock( io_requests_2_8_releaseLock ),
       .io_requests_8_grant( RRArbiter_2_io_requests_8_grant ),
       .io_requests_8_request( io_requests_2_8_request ),
       .io_requests_8_priorityLevel( io_requests_2_8_priorityLevel ),
       .io_requests_7_releaseLock( io_requests_2_7_releaseLock ),
       .io_requests_7_grant( RRArbiter_2_io_requests_7_grant ),
       .io_requests_7_request( io_requests_2_7_request ),
       .io_requests_7_priorityLevel( io_requests_2_7_priorityLevel ),
       .io_requests_6_releaseLock( io_requests_2_6_releaseLock ),
       .io_requests_6_grant( RRArbiter_2_io_requests_6_grant ),
       .io_requests_6_request( io_requests_2_6_request ),
       .io_requests_6_priorityLevel( io_requests_2_6_priorityLevel ),
       .io_requests_5_releaseLock( io_requests_2_5_releaseLock ),
       .io_requests_5_grant( RRArbiter_2_io_requests_5_grant ),
       .io_requests_5_request( io_requests_2_5_request ),
       .io_requests_5_priorityLevel( io_requests_2_5_priorityLevel ),
       .io_requests_4_releaseLock( io_requests_2_4_releaseLock ),
       .io_requests_4_grant( RRArbiter_2_io_requests_4_grant ),
       .io_requests_4_request( io_requests_2_4_request ),
       .io_requests_4_priorityLevel( io_requests_2_4_priorityLevel ),
       .io_requests_3_releaseLock( io_requests_2_3_releaseLock ),
       .io_requests_3_grant( RRArbiter_2_io_requests_3_grant ),
       .io_requests_3_request( io_requests_2_3_request ),
       .io_requests_3_priorityLevel( io_requests_2_3_priorityLevel ),
       .io_requests_2_releaseLock( io_requests_2_2_releaseLock ),
       .io_requests_2_grant( RRArbiter_2_io_requests_2_grant ),
       .io_requests_2_request( io_requests_2_2_request ),
       .io_requests_2_priorityLevel( io_requests_2_2_priorityLevel ),
       .io_requests_1_releaseLock( io_requests_2_1_releaseLock ),
       .io_requests_1_grant( RRArbiter_2_io_requests_1_grant ),
       .io_requests_1_request( io_requests_2_1_request ),
       .io_requests_1_priorityLevel( io_requests_2_1_priorityLevel ),
       .io_requests_0_releaseLock( io_requests_2_0_releaseLock ),
       .io_requests_0_grant( RRArbiter_2_io_requests_0_grant ),
       .io_requests_0_request( io_requests_2_0_request ),
       .io_requests_0_priorityLevel( io_requests_2_0_priorityLevel ),
       .io_resource_ready( io_resources_2_ready ),
       .io_resource_valid( RRArbiter_2_io_resource_valid ),
       .io_chosen( RRArbiter_2_io_chosen )
  );
  RRArbiter_1 RRArbiter_3(.clk(clk), .reset(reset),
       .io_requests_9_releaseLock( io_requests_3_9_releaseLock ),
       .io_requests_9_grant( RRArbiter_3_io_requests_9_grant ),
       .io_requests_9_request( io_requests_3_9_request ),
       .io_requests_9_priorityLevel( io_requests_3_9_priorityLevel ),
       .io_requests_8_releaseLock( io_requests_3_8_releaseLock ),
       .io_requests_8_grant( RRArbiter_3_io_requests_8_grant ),
       .io_requests_8_request( io_requests_3_8_request ),
       .io_requests_8_priorityLevel( io_requests_3_8_priorityLevel ),
       .io_requests_7_releaseLock( io_requests_3_7_releaseLock ),
       .io_requests_7_grant( RRArbiter_3_io_requests_7_grant ),
       .io_requests_7_request( io_requests_3_7_request ),
       .io_requests_7_priorityLevel( io_requests_3_7_priorityLevel ),
       .io_requests_6_releaseLock( io_requests_3_6_releaseLock ),
       .io_requests_6_grant( RRArbiter_3_io_requests_6_grant ),
       .io_requests_6_request( io_requests_3_6_request ),
       .io_requests_6_priorityLevel( io_requests_3_6_priorityLevel ),
       .io_requests_5_releaseLock( io_requests_3_5_releaseLock ),
       .io_requests_5_grant( RRArbiter_3_io_requests_5_grant ),
       .io_requests_5_request( io_requests_3_5_request ),
       .io_requests_5_priorityLevel( io_requests_3_5_priorityLevel ),
       .io_requests_4_releaseLock( io_requests_3_4_releaseLock ),
       .io_requests_4_grant( RRArbiter_3_io_requests_4_grant ),
       .io_requests_4_request( io_requests_3_4_request ),
       .io_requests_4_priorityLevel( io_requests_3_4_priorityLevel ),
       .io_requests_3_releaseLock( io_requests_3_3_releaseLock ),
       .io_requests_3_grant( RRArbiter_3_io_requests_3_grant ),
       .io_requests_3_request( io_requests_3_3_request ),
       .io_requests_3_priorityLevel( io_requests_3_3_priorityLevel ),
       .io_requests_2_releaseLock( io_requests_3_2_releaseLock ),
       .io_requests_2_grant( RRArbiter_3_io_requests_2_grant ),
       .io_requests_2_request( io_requests_3_2_request ),
       .io_requests_2_priorityLevel( io_requests_3_2_priorityLevel ),
       .io_requests_1_releaseLock( io_requests_3_1_releaseLock ),
       .io_requests_1_grant( RRArbiter_3_io_requests_1_grant ),
       .io_requests_1_request( io_requests_3_1_request ),
       .io_requests_1_priorityLevel( io_requests_3_1_priorityLevel ),
       .io_requests_0_releaseLock( io_requests_3_0_releaseLock ),
       .io_requests_0_grant( RRArbiter_3_io_requests_0_grant ),
       .io_requests_0_request( io_requests_3_0_request ),
       .io_requests_0_priorityLevel( io_requests_3_0_priorityLevel ),
       .io_resource_ready( io_resources_3_ready ),
       .io_resource_valid( RRArbiter_3_io_resource_valid ),
       .io_chosen( RRArbiter_3_io_chosen )
  );
  RRArbiter_1 RRArbiter_4(.clk(clk), .reset(reset),
       .io_requests_9_releaseLock( io_requests_4_9_releaseLock ),
       .io_requests_9_grant( RRArbiter_4_io_requests_9_grant ),
       .io_requests_9_request( io_requests_4_9_request ),
       .io_requests_9_priorityLevel( io_requests_4_9_priorityLevel ),
       .io_requests_8_releaseLock( io_requests_4_8_releaseLock ),
       .io_requests_8_grant( RRArbiter_4_io_requests_8_grant ),
       .io_requests_8_request( io_requests_4_8_request ),
       .io_requests_8_priorityLevel( io_requests_4_8_priorityLevel ),
       .io_requests_7_releaseLock( io_requests_4_7_releaseLock ),
       .io_requests_7_grant( RRArbiter_4_io_requests_7_grant ),
       .io_requests_7_request( io_requests_4_7_request ),
       .io_requests_7_priorityLevel( io_requests_4_7_priorityLevel ),
       .io_requests_6_releaseLock( io_requests_4_6_releaseLock ),
       .io_requests_6_grant( RRArbiter_4_io_requests_6_grant ),
       .io_requests_6_request( io_requests_4_6_request ),
       .io_requests_6_priorityLevel( io_requests_4_6_priorityLevel ),
       .io_requests_5_releaseLock( io_requests_4_5_releaseLock ),
       .io_requests_5_grant( RRArbiter_4_io_requests_5_grant ),
       .io_requests_5_request( io_requests_4_5_request ),
       .io_requests_5_priorityLevel( io_requests_4_5_priorityLevel ),
       .io_requests_4_releaseLock( io_requests_4_4_releaseLock ),
       .io_requests_4_grant( RRArbiter_4_io_requests_4_grant ),
       .io_requests_4_request( io_requests_4_4_request ),
       .io_requests_4_priorityLevel( io_requests_4_4_priorityLevel ),
       .io_requests_3_releaseLock( io_requests_4_3_releaseLock ),
       .io_requests_3_grant( RRArbiter_4_io_requests_3_grant ),
       .io_requests_3_request( io_requests_4_3_request ),
       .io_requests_3_priorityLevel( io_requests_4_3_priorityLevel ),
       .io_requests_2_releaseLock( io_requests_4_2_releaseLock ),
       .io_requests_2_grant( RRArbiter_4_io_requests_2_grant ),
       .io_requests_2_request( io_requests_4_2_request ),
       .io_requests_2_priorityLevel( io_requests_4_2_priorityLevel ),
       .io_requests_1_releaseLock( io_requests_4_1_releaseLock ),
       .io_requests_1_grant( RRArbiter_4_io_requests_1_grant ),
       .io_requests_1_request( io_requests_4_1_request ),
       .io_requests_1_priorityLevel( io_requests_4_1_priorityLevel ),
       .io_requests_0_releaseLock( io_requests_4_0_releaseLock ),
       .io_requests_0_grant( RRArbiter_4_io_requests_0_grant ),
       .io_requests_0_request( io_requests_4_0_request ),
       .io_requests_0_priorityLevel( io_requests_4_0_priorityLevel ),
       .io_resource_ready( io_resources_4_ready ),
       .io_resource_valid( RRArbiter_4_io_resource_valid ),
       .io_chosen( RRArbiter_4_io_chosen )
  );
  RRArbiter_1 RRArbiter_5(.clk(clk), .reset(reset),
       .io_requests_9_releaseLock( io_requests_5_9_releaseLock ),
       .io_requests_9_grant( RRArbiter_5_io_requests_9_grant ),
       .io_requests_9_request( io_requests_5_9_request ),
       .io_requests_9_priorityLevel( io_requests_5_9_priorityLevel ),
       .io_requests_8_releaseLock( io_requests_5_8_releaseLock ),
       .io_requests_8_grant( RRArbiter_5_io_requests_8_grant ),
       .io_requests_8_request( io_requests_5_8_request ),
       .io_requests_8_priorityLevel( io_requests_5_8_priorityLevel ),
       .io_requests_7_releaseLock( io_requests_5_7_releaseLock ),
       .io_requests_7_grant( RRArbiter_5_io_requests_7_grant ),
       .io_requests_7_request( io_requests_5_7_request ),
       .io_requests_7_priorityLevel( io_requests_5_7_priorityLevel ),
       .io_requests_6_releaseLock( io_requests_5_6_releaseLock ),
       .io_requests_6_grant( RRArbiter_5_io_requests_6_grant ),
       .io_requests_6_request( io_requests_5_6_request ),
       .io_requests_6_priorityLevel( io_requests_5_6_priorityLevel ),
       .io_requests_5_releaseLock( io_requests_5_5_releaseLock ),
       .io_requests_5_grant( RRArbiter_5_io_requests_5_grant ),
       .io_requests_5_request( io_requests_5_5_request ),
       .io_requests_5_priorityLevel( io_requests_5_5_priorityLevel ),
       .io_requests_4_releaseLock( io_requests_5_4_releaseLock ),
       .io_requests_4_grant( RRArbiter_5_io_requests_4_grant ),
       .io_requests_4_request( io_requests_5_4_request ),
       .io_requests_4_priorityLevel( io_requests_5_4_priorityLevel ),
       .io_requests_3_releaseLock( io_requests_5_3_releaseLock ),
       .io_requests_3_grant( RRArbiter_5_io_requests_3_grant ),
       .io_requests_3_request( io_requests_5_3_request ),
       .io_requests_3_priorityLevel( io_requests_5_3_priorityLevel ),
       .io_requests_2_releaseLock( io_requests_5_2_releaseLock ),
       .io_requests_2_grant( RRArbiter_5_io_requests_2_grant ),
       .io_requests_2_request( io_requests_5_2_request ),
       .io_requests_2_priorityLevel( io_requests_5_2_priorityLevel ),
       .io_requests_1_releaseLock( io_requests_5_1_releaseLock ),
       .io_requests_1_grant( RRArbiter_5_io_requests_1_grant ),
       .io_requests_1_request( io_requests_5_1_request ),
       .io_requests_1_priorityLevel( io_requests_5_1_priorityLevel ),
       .io_requests_0_releaseLock( io_requests_5_0_releaseLock ),
       .io_requests_0_grant( RRArbiter_5_io_requests_0_grant ),
       .io_requests_0_request( io_requests_5_0_request ),
       .io_requests_0_priorityLevel( io_requests_5_0_priorityLevel ),
       .io_resource_ready( io_resources_5_ready ),
       .io_resource_valid( RRArbiter_5_io_resource_valid ),
       .io_chosen( RRArbiter_5_io_chosen )
  );
  RRArbiter_1 RRArbiter_6(.clk(clk), .reset(reset),
       .io_requests_9_releaseLock( io_requests_6_9_releaseLock ),
       .io_requests_9_grant( RRArbiter_6_io_requests_9_grant ),
       .io_requests_9_request( io_requests_6_9_request ),
       .io_requests_9_priorityLevel( io_requests_6_9_priorityLevel ),
       .io_requests_8_releaseLock( io_requests_6_8_releaseLock ),
       .io_requests_8_grant( RRArbiter_6_io_requests_8_grant ),
       .io_requests_8_request( io_requests_6_8_request ),
       .io_requests_8_priorityLevel( io_requests_6_8_priorityLevel ),
       .io_requests_7_releaseLock( io_requests_6_7_releaseLock ),
       .io_requests_7_grant( RRArbiter_6_io_requests_7_grant ),
       .io_requests_7_request( io_requests_6_7_request ),
       .io_requests_7_priorityLevel( io_requests_6_7_priorityLevel ),
       .io_requests_6_releaseLock( io_requests_6_6_releaseLock ),
       .io_requests_6_grant( RRArbiter_6_io_requests_6_grant ),
       .io_requests_6_request( io_requests_6_6_request ),
       .io_requests_6_priorityLevel( io_requests_6_6_priorityLevel ),
       .io_requests_5_releaseLock( io_requests_6_5_releaseLock ),
       .io_requests_5_grant( RRArbiter_6_io_requests_5_grant ),
       .io_requests_5_request( io_requests_6_5_request ),
       .io_requests_5_priorityLevel( io_requests_6_5_priorityLevel ),
       .io_requests_4_releaseLock( io_requests_6_4_releaseLock ),
       .io_requests_4_grant( RRArbiter_6_io_requests_4_grant ),
       .io_requests_4_request( io_requests_6_4_request ),
       .io_requests_4_priorityLevel( io_requests_6_4_priorityLevel ),
       .io_requests_3_releaseLock( io_requests_6_3_releaseLock ),
       .io_requests_3_grant( RRArbiter_6_io_requests_3_grant ),
       .io_requests_3_request( io_requests_6_3_request ),
       .io_requests_3_priorityLevel( io_requests_6_3_priorityLevel ),
       .io_requests_2_releaseLock( io_requests_6_2_releaseLock ),
       .io_requests_2_grant( RRArbiter_6_io_requests_2_grant ),
       .io_requests_2_request( io_requests_6_2_request ),
       .io_requests_2_priorityLevel( io_requests_6_2_priorityLevel ),
       .io_requests_1_releaseLock( io_requests_6_1_releaseLock ),
       .io_requests_1_grant( RRArbiter_6_io_requests_1_grant ),
       .io_requests_1_request( io_requests_6_1_request ),
       .io_requests_1_priorityLevel( io_requests_6_1_priorityLevel ),
       .io_requests_0_releaseLock( io_requests_6_0_releaseLock ),
       .io_requests_0_grant( RRArbiter_6_io_requests_0_grant ),
       .io_requests_0_request( io_requests_6_0_request ),
       .io_requests_0_priorityLevel( io_requests_6_0_priorityLevel ),
       .io_resource_ready( io_resources_6_ready ),
       .io_resource_valid( RRArbiter_6_io_resource_valid ),
       .io_chosen( RRArbiter_6_io_chosen )
  );
  RRArbiter_1 RRArbiter_7(.clk(clk), .reset(reset),
       .io_requests_9_releaseLock( io_requests_7_9_releaseLock ),
       .io_requests_9_grant( RRArbiter_7_io_requests_9_grant ),
       .io_requests_9_request( io_requests_7_9_request ),
       .io_requests_9_priorityLevel( io_requests_7_9_priorityLevel ),
       .io_requests_8_releaseLock( io_requests_7_8_releaseLock ),
       .io_requests_8_grant( RRArbiter_7_io_requests_8_grant ),
       .io_requests_8_request( io_requests_7_8_request ),
       .io_requests_8_priorityLevel( io_requests_7_8_priorityLevel ),
       .io_requests_7_releaseLock( io_requests_7_7_releaseLock ),
       .io_requests_7_grant( RRArbiter_7_io_requests_7_grant ),
       .io_requests_7_request( io_requests_7_7_request ),
       .io_requests_7_priorityLevel( io_requests_7_7_priorityLevel ),
       .io_requests_6_releaseLock( io_requests_7_6_releaseLock ),
       .io_requests_6_grant( RRArbiter_7_io_requests_6_grant ),
       .io_requests_6_request( io_requests_7_6_request ),
       .io_requests_6_priorityLevel( io_requests_7_6_priorityLevel ),
       .io_requests_5_releaseLock( io_requests_7_5_releaseLock ),
       .io_requests_5_grant( RRArbiter_7_io_requests_5_grant ),
       .io_requests_5_request( io_requests_7_5_request ),
       .io_requests_5_priorityLevel( io_requests_7_5_priorityLevel ),
       .io_requests_4_releaseLock( io_requests_7_4_releaseLock ),
       .io_requests_4_grant( RRArbiter_7_io_requests_4_grant ),
       .io_requests_4_request( io_requests_7_4_request ),
       .io_requests_4_priorityLevel( io_requests_7_4_priorityLevel ),
       .io_requests_3_releaseLock( io_requests_7_3_releaseLock ),
       .io_requests_3_grant( RRArbiter_7_io_requests_3_grant ),
       .io_requests_3_request( io_requests_7_3_request ),
       .io_requests_3_priorityLevel( io_requests_7_3_priorityLevel ),
       .io_requests_2_releaseLock( io_requests_7_2_releaseLock ),
       .io_requests_2_grant( RRArbiter_7_io_requests_2_grant ),
       .io_requests_2_request( io_requests_7_2_request ),
       .io_requests_2_priorityLevel( io_requests_7_2_priorityLevel ),
       .io_requests_1_releaseLock( io_requests_7_1_releaseLock ),
       .io_requests_1_grant( RRArbiter_7_io_requests_1_grant ),
       .io_requests_1_request( io_requests_7_1_request ),
       .io_requests_1_priorityLevel( io_requests_7_1_priorityLevel ),
       .io_requests_0_releaseLock( io_requests_7_0_releaseLock ),
       .io_requests_0_grant( RRArbiter_7_io_requests_0_grant ),
       .io_requests_0_request( io_requests_7_0_request ),
       .io_requests_0_priorityLevel( io_requests_7_0_priorityLevel ),
       .io_resource_ready( io_resources_7_ready ),
       .io_resource_valid( RRArbiter_7_io_resource_valid ),
       .io_chosen( RRArbiter_7_io_chosen )
  );
  RRArbiter_1 RRArbiter_8(.clk(clk), .reset(reset),
       .io_requests_9_releaseLock( io_requests_8_9_releaseLock ),
       .io_requests_9_grant( RRArbiter_8_io_requests_9_grant ),
       .io_requests_9_request( io_requests_8_9_request ),
       .io_requests_9_priorityLevel( io_requests_8_9_priorityLevel ),
       .io_requests_8_releaseLock( io_requests_8_8_releaseLock ),
       .io_requests_8_grant( RRArbiter_8_io_requests_8_grant ),
       .io_requests_8_request( io_requests_8_8_request ),
       .io_requests_8_priorityLevel( io_requests_8_8_priorityLevel ),
       .io_requests_7_releaseLock( io_requests_8_7_releaseLock ),
       .io_requests_7_grant( RRArbiter_8_io_requests_7_grant ),
       .io_requests_7_request( io_requests_8_7_request ),
       .io_requests_7_priorityLevel( io_requests_8_7_priorityLevel ),
       .io_requests_6_releaseLock( io_requests_8_6_releaseLock ),
       .io_requests_6_grant( RRArbiter_8_io_requests_6_grant ),
       .io_requests_6_request( io_requests_8_6_request ),
       .io_requests_6_priorityLevel( io_requests_8_6_priorityLevel ),
       .io_requests_5_releaseLock( io_requests_8_5_releaseLock ),
       .io_requests_5_grant( RRArbiter_8_io_requests_5_grant ),
       .io_requests_5_request( io_requests_8_5_request ),
       .io_requests_5_priorityLevel( io_requests_8_5_priorityLevel ),
       .io_requests_4_releaseLock( io_requests_8_4_releaseLock ),
       .io_requests_4_grant( RRArbiter_8_io_requests_4_grant ),
       .io_requests_4_request( io_requests_8_4_request ),
       .io_requests_4_priorityLevel( io_requests_8_4_priorityLevel ),
       .io_requests_3_releaseLock( io_requests_8_3_releaseLock ),
       .io_requests_3_grant( RRArbiter_8_io_requests_3_grant ),
       .io_requests_3_request( io_requests_8_3_request ),
       .io_requests_3_priorityLevel( io_requests_8_3_priorityLevel ),
       .io_requests_2_releaseLock( io_requests_8_2_releaseLock ),
       .io_requests_2_grant( RRArbiter_8_io_requests_2_grant ),
       .io_requests_2_request( io_requests_8_2_request ),
       .io_requests_2_priorityLevel( io_requests_8_2_priorityLevel ),
       .io_requests_1_releaseLock( io_requests_8_1_releaseLock ),
       .io_requests_1_grant( RRArbiter_8_io_requests_1_grant ),
       .io_requests_1_request( io_requests_8_1_request ),
       .io_requests_1_priorityLevel( io_requests_8_1_priorityLevel ),
       .io_requests_0_releaseLock( io_requests_8_0_releaseLock ),
       .io_requests_0_grant( RRArbiter_8_io_requests_0_grant ),
       .io_requests_0_request( io_requests_8_0_request ),
       .io_requests_0_priorityLevel( io_requests_8_0_priorityLevel ),
       .io_resource_ready( io_resources_8_ready ),
       .io_resource_valid( RRArbiter_8_io_resource_valid ),
       .io_chosen( RRArbiter_8_io_chosen )
  );
  RRArbiter_1 RRArbiter_9(.clk(clk), .reset(reset),
       .io_requests_9_releaseLock( io_requests_9_9_releaseLock ),
       .io_requests_9_grant( RRArbiter_9_io_requests_9_grant ),
       .io_requests_9_request( io_requests_9_9_request ),
       .io_requests_9_priorityLevel( io_requests_9_9_priorityLevel ),
       .io_requests_8_releaseLock( io_requests_9_8_releaseLock ),
       .io_requests_8_grant( RRArbiter_9_io_requests_8_grant ),
       .io_requests_8_request( io_requests_9_8_request ),
       .io_requests_8_priorityLevel( io_requests_9_8_priorityLevel ),
       .io_requests_7_releaseLock( io_requests_9_7_releaseLock ),
       .io_requests_7_grant( RRArbiter_9_io_requests_7_grant ),
       .io_requests_7_request( io_requests_9_7_request ),
       .io_requests_7_priorityLevel( io_requests_9_7_priorityLevel ),
       .io_requests_6_releaseLock( io_requests_9_6_releaseLock ),
       .io_requests_6_grant( RRArbiter_9_io_requests_6_grant ),
       .io_requests_6_request( io_requests_9_6_request ),
       .io_requests_6_priorityLevel( io_requests_9_6_priorityLevel ),
       .io_requests_5_releaseLock( io_requests_9_5_releaseLock ),
       .io_requests_5_grant( RRArbiter_9_io_requests_5_grant ),
       .io_requests_5_request( io_requests_9_5_request ),
       .io_requests_5_priorityLevel( io_requests_9_5_priorityLevel ),
       .io_requests_4_releaseLock( io_requests_9_4_releaseLock ),
       .io_requests_4_grant( RRArbiter_9_io_requests_4_grant ),
       .io_requests_4_request( io_requests_9_4_request ),
       .io_requests_4_priorityLevel( io_requests_9_4_priorityLevel ),
       .io_requests_3_releaseLock( io_requests_9_3_releaseLock ),
       .io_requests_3_grant( RRArbiter_9_io_requests_3_grant ),
       .io_requests_3_request( io_requests_9_3_request ),
       .io_requests_3_priorityLevel( io_requests_9_3_priorityLevel ),
       .io_requests_2_releaseLock( io_requests_9_2_releaseLock ),
       .io_requests_2_grant( RRArbiter_9_io_requests_2_grant ),
       .io_requests_2_request( io_requests_9_2_request ),
       .io_requests_2_priorityLevel( io_requests_9_2_priorityLevel ),
       .io_requests_1_releaseLock( io_requests_9_1_releaseLock ),
       .io_requests_1_grant( RRArbiter_9_io_requests_1_grant ),
       .io_requests_1_request( io_requests_9_1_request ),
       .io_requests_1_priorityLevel( io_requests_9_1_priorityLevel ),
       .io_requests_0_releaseLock( io_requests_9_0_releaseLock ),
       .io_requests_0_grant( RRArbiter_9_io_requests_0_grant ),
       .io_requests_0_request( io_requests_9_0_request ),
       .io_requests_0_priorityLevel( io_requests_9_0_priorityLevel ),
       .io_resource_ready( io_resources_9_ready ),
       .io_resource_valid( RRArbiter_9_io_resource_valid ),
       .io_chosen( RRArbiter_9_io_chosen )
  );
endmodule

module VCRouterOutputStateManagement(input clk, input reset,
    input  io_swAllocGranted,
    input  io_creditsAvail,
    output[1:0] io_currentState
);

  reg [1:0] curState;
  wire[1:0] T36;
  wire[1:0] T0;
  wire[1:0] T1;
  wire[1:0] T2;
  wire[1:0] T3;
  wire[1:0] T4;
  wire[1:0] T5;
  wire[1:0] T6;
  wire[1:0] T7;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    curState = {1{1'b0}};
  end
// synthesis translate_on
`endif

  assign io_currentState = curState;
  assign T36 = reset ? 2'h0 : T0;
  assign T0 = T34 ? 2'h3 : T1;
  assign T1 = T29 ? 2'h2 : T2;
  assign T2 = T26 ? 2'h3 : T3;
  assign T3 = T22 ? 2'h0 : T4;
  assign T4 = T16 ? 2'h2 : T5;
  assign T5 = T13 ? 2'h2 : T6;
  assign T6 = T11 ? 2'h0 : T7;
  assign T7 = T8 ? 2'h1 : curState;
  assign T8 = T10 & T9;
  assign T9 = io_swAllocGranted & io_creditsAvail;
  assign T10 = curState == 2'h0;
  assign T11 = T10 & T12;
  assign T12 = T9 ^ 1'h1;
  assign T13 = T15 & T14;
  assign T14 = curState == 2'h1;
  assign T15 = T10 ^ 1'h1;
  assign T16 = T18 & T17;
  assign T17 = io_creditsAvail & io_swAllocGranted;
  assign T18 = T20 & T19;
  assign T19 = curState == 2'h2;
  assign T20 = T21 ^ 1'h1;
  assign T21 = T10 | T14;
  assign T22 = T18 & T23;
  assign T23 = T25 & T24;
  assign T24 = ~ io_swAllocGranted;
  assign T25 = T17 ^ 1'h1;
  assign T26 = T18 & T27;
  assign T27 = T28 ^ 1'h1;
  assign T28 = T17 | T24;
  assign T29 = T30 & io_creditsAvail;
  assign T30 = T32 & T31;
  assign T31 = curState == 2'h3;
  assign T32 = T33 ^ 1'h1;
  assign T33 = T21 | T19;
  assign T34 = T30 & T35;
  assign T35 = io_creditsAvail ^ 1'h1;

  always @(posedge clk) begin
    if(reset) begin
      curState <= 2'h0;
    end else if(T34) begin
      curState <= 2'h3;
    end else if(T29) begin
      curState <= 2'h2;
    end else if(T26) begin
      curState <= 2'h3;
    end else if(T22) begin
      curState <= 2'h0;
    end else if(T16) begin
      curState <= 2'h2;
    end else if(T13) begin
      curState <= 2'h2;
    end else if(T11) begin
      curState <= 2'h0;
    end else if(T8) begin
      curState <= 2'h1;
    end
  end
endmodule

module CreditGen(
    output io_outCredit_grant,
    input  io_inGrant
);



  assign io_outCredit_grant = io_inGrant;
endmodule

module RouterRegFile(input clk, input reset,
    input [54:0] io_writeData,
    input  io_writeEnable,
    output io_full,
    output[54:0] io_readData,
    output io_readValid,
    input  io_readIncrement,
    input [54:0] io_writePipelineReg_2,
    input [54:0] io_writePipelineReg_1,
    input [54:0] io_writePipelineReg_0,
    input  io_wePipelineReg_2,
    input  io_wePipelineReg_1,
    input  io_wePipelineReg_0,
    output[54:0] io_readPipelineReg_2,
    output[54:0] io_readPipelineReg_1,
    output[54:0] io_readPipelineReg_0,
    output io_rvPipelineReg_2,
    output io_rvPipelineReg_1,
    output io_rvPipelineReg_0
);

  reg  regRVPipelineRegs_0;
  reg  regRVPipelineRegs_1;
  reg  regRVPipelineRegs_2;
  reg [54:0] regPipelineRegs_0;
  wire[54:0] T244;
  reg [54:0] regPipelineRegs_1;
  wire[54:0] T245;
  reg [54:0] regPipelineRegs_2;
  wire[54:0] T246;
  wire T0;
  wire T1;
  wire[15:0] T2;
  wire[15:0] T3;
  wire[7:0] T4;
  wire[3:0] T5;
  wire[1:0] T6;
  reg  regFileValid_0;
  wire T247;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  wire[15:0] T11;
  wire[3:0] T12;
  reg [3:0] writePointer;
  wire[3:0] T248;
  wire[3:0] T13;
  wire[3:0] T14;
  wire[3:0] T15;
  wire T16;
  wire T17;
  wire[4:0] T249;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  reg  regFileValid_2;
  wire T250;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire[15:0] T32;
  wire[3:0] T33;
  reg [3:0] readPointer;
  wire[3:0] T251;
  wire[3:0] T34;
  wire[3:0] T35;
  wire[3:0] T36;
  wire T37;
  wire T38;
  wire[4:0] T252;
  reg  regFileValid_3;
  wire T253;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  reg  regFileValid_4;
  wire T254;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  reg  regFileValid_5;
  wire T255;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire T61;
  wire T62;
  reg  regFileValid_6;
  wire T256;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire T67;
  wire T68;
  reg  regFileValid_7;
  wire T257;
  wire T69;
  wire T70;
  wire T71;
  wire T72;
  wire T73;
  wire T74;
  wire T75;
  wire T76;
  wire T77;
  wire T78;
  wire T79;
  wire T80;
  reg  regFileValid_8;
  wire T258;
  wire T81;
  wire T82;
  wire T83;
  wire T84;
  wire T85;
  wire T86;
  reg  regFileValid_9;
  wire T259;
  wire T87;
  wire T88;
  wire T89;
  wire T90;
  wire T91;
  wire T92;
  wire T93;
  wire T94;
  reg  regFileValid_10;
  wire T260;
  wire T95;
  wire T96;
  wire T97;
  wire T98;
  wire T99;
  wire T100;
  reg  regFileValid_11;
  wire T261;
  wire T101;
  wire T102;
  wire T103;
  wire T104;
  wire T105;
  wire T106;
  wire T107;
  wire T108;
  wire T109;
  wire T110;
  reg  regFileValid_12;
  wire T262;
  wire T111;
  wire T112;
  wire T113;
  wire T114;
  wire T115;
  wire T116;
  reg  regFileValid_13;
  wire T263;
  wire T117;
  wire T118;
  wire T119;
  wire T120;
  wire T121;
  wire T122;
  wire T123;
  wire T124;
  reg  regFileValid_14;
  wire T264;
  wire T125;
  wire T126;
  wire T127;
  wire T128;
  wire T129;
  wire T130;
  reg  regFileValid_15;
  wire T265;
  wire T131;
  wire T132;
  wire T133;
  wire T134;
  wire T135;
  wire T136;
  wire T137;
  wire T138;
  wire T139;
  wire T140;
  wire T141;
  wire T142;
  reg  regFileValid_1;
  wire T266;
  wire T143;
  wire T144;
  wire T145;
  wire T146;
  wire T147;
  wire T148;
  wire[1:0] T149;
  wire[3:0] T150;
  wire[1:0] T151;
  wire[1:0] T152;
  wire[7:0] T153;
  wire[3:0] T154;
  wire[1:0] T155;
  wire[1:0] T156;
  wire[3:0] T157;
  wire[1:0] T158;
  wire[1:0] T159;
  wire T160;
  wire[54:0] T161;
  wire[54:0] T162;
  wire[54:0] T163;
  wire[54:0] T164;
  reg [54:0] regFile_0;
  wire[54:0] T267;
  wire[54:0] T165;
  wire T166;
  wire T167;
  wire[15:0] T168;
  wire[3:0] T169;
  reg [54:0] regFile_1;
  wire[54:0] T268;
  wire[54:0] T170;
  wire T171;
  wire T172;
  wire T173;
  wire[3:0] T174;
  wire[54:0] T175;
  reg [54:0] regFile_2;
  wire[54:0] T269;
  wire[54:0] T176;
  wire T177;
  wire T178;
  reg [54:0] regFile_3;
  wire[54:0] T270;
  wire[54:0] T179;
  wire T180;
  wire T181;
  wire T182;
  wire T183;
  wire[54:0] T184;
  wire[54:0] T185;
  reg [54:0] regFile_4;
  wire[54:0] T271;
  wire[54:0] T186;
  wire T187;
  wire T188;
  reg [54:0] regFile_5;
  wire[54:0] T272;
  wire[54:0] T189;
  wire T190;
  wire T191;
  wire T192;
  wire[54:0] T193;
  reg [54:0] regFile_6;
  wire[54:0] T273;
  wire[54:0] T194;
  wire T195;
  wire T196;
  reg [54:0] regFile_7;
  wire[54:0] T274;
  wire[54:0] T197;
  wire T198;
  wire T199;
  wire T200;
  wire T201;
  wire T202;
  wire[54:0] T203;
  wire[54:0] T204;
  wire[54:0] T205;
  reg [54:0] regFile_8;
  wire[54:0] T275;
  wire[54:0] T206;
  wire T207;
  wire T208;
  reg [54:0] regFile_9;
  wire[54:0] T276;
  wire[54:0] T209;
  wire T210;
  wire T211;
  wire T212;
  wire[54:0] T213;
  reg [54:0] regFile_10;
  wire[54:0] T277;
  wire[54:0] T214;
  wire T215;
  wire T216;
  reg [54:0] regFile_11;
  wire[54:0] T278;
  wire[54:0] T217;
  wire T218;
  wire T219;
  wire T220;
  wire T221;
  wire[54:0] T222;
  wire[54:0] T223;
  reg [54:0] regFile_12;
  wire[54:0] T279;
  wire[54:0] T224;
  wire T225;
  wire T226;
  reg [54:0] regFile_13;
  wire[54:0] T280;
  wire[54:0] T227;
  wire T228;
  wire T229;
  wire T230;
  wire[54:0] T231;
  reg [54:0] regFile_14;
  wire[54:0] T281;
  wire[54:0] T232;
  wire T233;
  wire T234;
  reg [54:0] regFile_15;
  wire[54:0] T282;
  wire[54:0] T235;
  wire T236;
  wire T237;
  wire T238;
  wire T239;
  wire T240;
  wire T241;
  wire T242;
  wire[15:0] T243;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    regRVPipelineRegs_0 = {1{1'b0}};
    regRVPipelineRegs_1 = {1{1'b0}};
    regRVPipelineRegs_2 = {1{1'b0}};
    regPipelineRegs_0 = {2{1'b0}};
    regPipelineRegs_1 = {2{1'b0}};
    regPipelineRegs_2 = {2{1'b0}};
    regFileValid_0 = {1{1'b0}};
    writePointer = {1{1'b0}};
    regFileValid_2 = {1{1'b0}};
    readPointer = {1{1'b0}};
    regFileValid_3 = {1{1'b0}};
    regFileValid_4 = {1{1'b0}};
    regFileValid_5 = {1{1'b0}};
    regFileValid_6 = {1{1'b0}};
    regFileValid_7 = {1{1'b0}};
    regFileValid_8 = {1{1'b0}};
    regFileValid_9 = {1{1'b0}};
    regFileValid_10 = {1{1'b0}};
    regFileValid_11 = {1{1'b0}};
    regFileValid_12 = {1{1'b0}};
    regFileValid_13 = {1{1'b0}};
    regFileValid_14 = {1{1'b0}};
    regFileValid_15 = {1{1'b0}};
    regFileValid_1 = {1{1'b0}};
    regFile_0 = {2{1'b0}};
    regFile_1 = {2{1'b0}};
    regFile_2 = {2{1'b0}};
    regFile_3 = {2{1'b0}};
    regFile_4 = {2{1'b0}};
    regFile_5 = {2{1'b0}};
    regFile_6 = {2{1'b0}};
    regFile_7 = {2{1'b0}};
    regFile_8 = {2{1'b0}};
    regFile_9 = {2{1'b0}};
    regFile_10 = {2{1'b0}};
    regFile_11 = {2{1'b0}};
    regFile_12 = {2{1'b0}};
    regFile_13 = {2{1'b0}};
    regFile_14 = {2{1'b0}};
    regFile_15 = {2{1'b0}};
  end
// synthesis translate_on
`endif

  assign io_rvPipelineReg_0 = regRVPipelineRegs_0;
  assign io_rvPipelineReg_1 = regRVPipelineRegs_1;
  assign io_rvPipelineReg_2 = regRVPipelineRegs_2;
  assign io_readPipelineReg_0 = regPipelineRegs_0;
  assign T244 = reset ? 55'h0 : io_writePipelineReg_0;
  assign io_readPipelineReg_1 = regPipelineRegs_1;
  assign T245 = reset ? 55'h0 : io_writePipelineReg_1;
  assign io_readPipelineReg_2 = regPipelineRegs_2;
  assign T246 = reset ? 55'h0 : io_writePipelineReg_2;
  assign io_readValid = T0;
  assign T0 = T160 & T1;
  assign T1 = T2 != 16'h0;
  assign T2 = T3;
  assign T3 = {T153, T4};
  assign T4 = {T150, T5};
  assign T5 = {T149, T6};
  assign T6 = {regFileValid_1, regFileValid_0};
  assign T247 = reset ? 1'h0 : T7;
  assign T7 = T141 ? 1'h0 : T8;
  assign T8 = T9 ? 1'h1 : regFileValid_0;
  assign T9 = T18 & T10;
  assign T10 = T11[1'h0:1'h0];
  assign T11 = 1'h1 << T12;
  assign T12 = writePointer;
  assign T248 = reset ? 4'h0 : T13;
  assign T13 = T16 ? 4'h0 : T14;
  assign T14 = T18 ? T15 : writePointer;
  assign T15 = writePointer + 4'h1;
  assign T16 = T18 & T17;
  assign T17 = T249 == 5'h10;
  assign T249 = {1'h0, writePointer};
  assign T18 = io_writeEnable & T19;
  assign T19 = T20 ^ 1'h1;
  assign T20 = T140 ? T78 : T21;
  assign T21 = T77 ? T47 : T22;
  assign T22 = T46 ? T25 : T23;
  assign T23 = T24 ? regFileValid_1 : regFileValid_0;
  assign T24 = T12[1'h0:1'h0];
  assign T25 = T45 ? regFileValid_3 : regFileValid_2;
  assign T250 = reset ? 1'h0 : T26;
  assign T26 = T30 ? 1'h0 : T27;
  assign T27 = T28 ? 1'h1 : regFileValid_2;
  assign T28 = T18 & T29;
  assign T29 = T11[2'h2:2'h2];
  assign T30 = io_readIncrement & T31;
  assign T31 = T32[2'h2:2'h2];
  assign T32 = 1'h1 << T33;
  assign T33 = readPointer;
  assign T251 = reset ? 4'h0 : T34;
  assign T34 = T37 ? 4'h0 : T35;
  assign T35 = io_readIncrement ? T36 : readPointer;
  assign T36 = readPointer + 4'h1;
  assign T37 = io_readIncrement & T38;
  assign T38 = T252 == 5'h10;
  assign T252 = {1'h0, readPointer};
  assign T253 = reset ? 1'h0 : T39;
  assign T39 = T43 ? 1'h0 : T40;
  assign T40 = T41 ? 1'h1 : regFileValid_3;
  assign T41 = T18 & T42;
  assign T42 = T11[2'h3:2'h3];
  assign T43 = io_readIncrement & T44;
  assign T44 = T32[2'h3:2'h3];
  assign T45 = T12[1'h0:1'h0];
  assign T46 = T12[1'h1:1'h1];
  assign T47 = T76 ? T62 : T48;
  assign T48 = T61 ? regFileValid_5 : regFileValid_4;
  assign T254 = reset ? 1'h0 : T49;
  assign T49 = T53 ? 1'h0 : T50;
  assign T50 = T51 ? 1'h1 : regFileValid_4;
  assign T51 = T18 & T52;
  assign T52 = T11[3'h4:3'h4];
  assign T53 = io_readIncrement & T54;
  assign T54 = T32[3'h4:3'h4];
  assign T255 = reset ? 1'h0 : T55;
  assign T55 = T59 ? 1'h0 : T56;
  assign T56 = T57 ? 1'h1 : regFileValid_5;
  assign T57 = T18 & T58;
  assign T58 = T11[3'h5:3'h5];
  assign T59 = io_readIncrement & T60;
  assign T60 = T32[3'h5:3'h5];
  assign T61 = T12[1'h0:1'h0];
  assign T62 = T75 ? regFileValid_7 : regFileValid_6;
  assign T256 = reset ? 1'h0 : T63;
  assign T63 = T67 ? 1'h0 : T64;
  assign T64 = T65 ? 1'h1 : regFileValid_6;
  assign T65 = T18 & T66;
  assign T66 = T11[3'h6:3'h6];
  assign T67 = io_readIncrement & T68;
  assign T68 = T32[3'h6:3'h6];
  assign T257 = reset ? 1'h0 : T69;
  assign T69 = T73 ? 1'h0 : T70;
  assign T70 = T71 ? 1'h1 : regFileValid_7;
  assign T71 = T18 & T72;
  assign T72 = T11[3'h7:3'h7];
  assign T73 = io_readIncrement & T74;
  assign T74 = T32[3'h7:3'h7];
  assign T75 = T12[1'h0:1'h0];
  assign T76 = T12[1'h1:1'h1];
  assign T77 = T12[2'h2:2'h2];
  assign T78 = T139 ? T109 : T79;
  assign T79 = T108 ? T94 : T80;
  assign T80 = T93 ? regFileValid_9 : regFileValid_8;
  assign T258 = reset ? 1'h0 : T81;
  assign T81 = T85 ? 1'h0 : T82;
  assign T82 = T83 ? 1'h1 : regFileValid_8;
  assign T83 = T18 & T84;
  assign T84 = T11[4'h8:4'h8];
  assign T85 = io_readIncrement & T86;
  assign T86 = T32[4'h8:4'h8];
  assign T259 = reset ? 1'h0 : T87;
  assign T87 = T91 ? 1'h0 : T88;
  assign T88 = T89 ? 1'h1 : regFileValid_9;
  assign T89 = T18 & T90;
  assign T90 = T11[4'h9:4'h9];
  assign T91 = io_readIncrement & T92;
  assign T92 = T32[4'h9:4'h9];
  assign T93 = T12[1'h0:1'h0];
  assign T94 = T107 ? regFileValid_11 : regFileValid_10;
  assign T260 = reset ? 1'h0 : T95;
  assign T95 = T99 ? 1'h0 : T96;
  assign T96 = T97 ? 1'h1 : regFileValid_10;
  assign T97 = T18 & T98;
  assign T98 = T11[4'ha:4'ha];
  assign T99 = io_readIncrement & T100;
  assign T100 = T32[4'ha:4'ha];
  assign T261 = reset ? 1'h0 : T101;
  assign T101 = T105 ? 1'h0 : T102;
  assign T102 = T103 ? 1'h1 : regFileValid_11;
  assign T103 = T18 & T104;
  assign T104 = T11[4'hb:4'hb];
  assign T105 = io_readIncrement & T106;
  assign T106 = T32[4'hb:4'hb];
  assign T107 = T12[1'h0:1'h0];
  assign T108 = T12[1'h1:1'h1];
  assign T109 = T138 ? T124 : T110;
  assign T110 = T123 ? regFileValid_13 : regFileValid_12;
  assign T262 = reset ? 1'h0 : T111;
  assign T111 = T115 ? 1'h0 : T112;
  assign T112 = T113 ? 1'h1 : regFileValid_12;
  assign T113 = T18 & T114;
  assign T114 = T11[4'hc:4'hc];
  assign T115 = io_readIncrement & T116;
  assign T116 = T32[4'hc:4'hc];
  assign T263 = reset ? 1'h0 : T117;
  assign T117 = T121 ? 1'h0 : T118;
  assign T118 = T119 ? 1'h1 : regFileValid_13;
  assign T119 = T18 & T120;
  assign T120 = T11[4'hd:4'hd];
  assign T121 = io_readIncrement & T122;
  assign T122 = T32[4'hd:4'hd];
  assign T123 = T12[1'h0:1'h0];
  assign T124 = T137 ? regFileValid_15 : regFileValid_14;
  assign T264 = reset ? 1'h0 : T125;
  assign T125 = T129 ? 1'h0 : T126;
  assign T126 = T127 ? 1'h1 : regFileValid_14;
  assign T127 = T18 & T128;
  assign T128 = T11[4'he:4'he];
  assign T129 = io_readIncrement & T130;
  assign T130 = T32[4'he:4'he];
  assign T265 = reset ? 1'h0 : T131;
  assign T131 = T135 ? 1'h0 : T132;
  assign T132 = T133 ? 1'h1 : regFileValid_15;
  assign T133 = T18 & T134;
  assign T134 = T11[4'hf:4'hf];
  assign T135 = io_readIncrement & T136;
  assign T136 = T32[4'hf:4'hf];
  assign T137 = T12[1'h0:1'h0];
  assign T138 = T12[1'h1:1'h1];
  assign T139 = T12[2'h2:2'h2];
  assign T140 = T12[2'h3:2'h3];
  assign T141 = io_readIncrement & T142;
  assign T142 = T32[1'h0:1'h0];
  assign T266 = reset ? 1'h0 : T143;
  assign T143 = T147 ? 1'h0 : T144;
  assign T144 = T145 ? 1'h1 : regFileValid_1;
  assign T145 = T18 & T146;
  assign T146 = T11[1'h1:1'h1];
  assign T147 = io_readIncrement & T148;
  assign T148 = T32[1'h1:1'h1];
  assign T149 = {regFileValid_3, regFileValid_2};
  assign T150 = {T152, T151};
  assign T151 = {regFileValid_5, regFileValid_4};
  assign T152 = {regFileValid_7, regFileValid_6};
  assign T153 = {T157, T154};
  assign T154 = {T156, T155};
  assign T155 = {regFileValid_9, regFileValid_8};
  assign T156 = {regFileValid_11, regFileValid_10};
  assign T157 = {T159, T158};
  assign T158 = {regFileValid_13, regFileValid_12};
  assign T159 = {regFileValid_15, regFileValid_14};
  assign T160 = writePointer != readPointer;
  assign io_readData = T161;
  assign T161 = T241 ? T203 : T162;
  assign T162 = T202 ? T184 : T163;
  assign T163 = T183 ? T175 : T164;
  assign T164 = T173 ? regFile_1 : regFile_0;
  assign T267 = reset ? 55'h0 : T165;
  assign T165 = T166 ? io_writeData : regFile_0;
  assign T166 = T18 & T167;
  assign T167 = T168[1'h0:1'h0];
  assign T168 = 1'h1 << T169;
  assign T169 = writePointer;
  assign T268 = reset ? 55'h0 : T170;
  assign T170 = T171 ? io_writeData : regFile_1;
  assign T171 = T18 & T172;
  assign T172 = T168[1'h1:1'h1];
  assign T173 = T174[1'h0:1'h0];
  assign T174 = readPointer;
  assign T175 = T182 ? regFile_3 : regFile_2;
  assign T269 = reset ? 55'h0 : T176;
  assign T176 = T177 ? io_writeData : regFile_2;
  assign T177 = T18 & T178;
  assign T178 = T168[2'h2:2'h2];
  assign T270 = reset ? 55'h0 : T179;
  assign T179 = T180 ? io_writeData : regFile_3;
  assign T180 = T18 & T181;
  assign T181 = T168[2'h3:2'h3];
  assign T182 = T174[1'h0:1'h0];
  assign T183 = T174[1'h1:1'h1];
  assign T184 = T201 ? T193 : T185;
  assign T185 = T192 ? regFile_5 : regFile_4;
  assign T271 = reset ? 55'h0 : T186;
  assign T186 = T187 ? io_writeData : regFile_4;
  assign T187 = T18 & T188;
  assign T188 = T168[3'h4:3'h4];
  assign T272 = reset ? 55'h0 : T189;
  assign T189 = T190 ? io_writeData : regFile_5;
  assign T190 = T18 & T191;
  assign T191 = T168[3'h5:3'h5];
  assign T192 = T174[1'h0:1'h0];
  assign T193 = T200 ? regFile_7 : regFile_6;
  assign T273 = reset ? 55'h0 : T194;
  assign T194 = T195 ? io_writeData : regFile_6;
  assign T195 = T18 & T196;
  assign T196 = T168[3'h6:3'h6];
  assign T274 = reset ? 55'h0 : T197;
  assign T197 = T198 ? io_writeData : regFile_7;
  assign T198 = T18 & T199;
  assign T199 = T168[3'h7:3'h7];
  assign T200 = T174[1'h0:1'h0];
  assign T201 = T174[1'h1:1'h1];
  assign T202 = T174[2'h2:2'h2];
  assign T203 = T240 ? T222 : T204;
  assign T204 = T221 ? T213 : T205;
  assign T205 = T212 ? regFile_9 : regFile_8;
  assign T275 = reset ? 55'h0 : T206;
  assign T206 = T207 ? io_writeData : regFile_8;
  assign T207 = T18 & T208;
  assign T208 = T168[4'h8:4'h8];
  assign T276 = reset ? 55'h0 : T209;
  assign T209 = T210 ? io_writeData : regFile_9;
  assign T210 = T18 & T211;
  assign T211 = T168[4'h9:4'h9];
  assign T212 = T174[1'h0:1'h0];
  assign T213 = T220 ? regFile_11 : regFile_10;
  assign T277 = reset ? 55'h0 : T214;
  assign T214 = T215 ? io_writeData : regFile_10;
  assign T215 = T18 & T216;
  assign T216 = T168[4'ha:4'ha];
  assign T278 = reset ? 55'h0 : T217;
  assign T217 = T218 ? io_writeData : regFile_11;
  assign T218 = T18 & T219;
  assign T219 = T168[4'hb:4'hb];
  assign T220 = T174[1'h0:1'h0];
  assign T221 = T174[1'h1:1'h1];
  assign T222 = T239 ? T231 : T223;
  assign T223 = T230 ? regFile_13 : regFile_12;
  assign T279 = reset ? 55'h0 : T224;
  assign T224 = T225 ? io_writeData : regFile_12;
  assign T225 = T18 & T226;
  assign T226 = T168[4'hc:4'hc];
  assign T280 = reset ? 55'h0 : T227;
  assign T227 = T228 ? io_writeData : regFile_13;
  assign T228 = T18 & T229;
  assign T229 = T168[4'hd:4'hd];
  assign T230 = T174[1'h0:1'h0];
  assign T231 = T238 ? regFile_15 : regFile_14;
  assign T281 = reset ? 55'h0 : T232;
  assign T232 = T233 ? io_writeData : regFile_14;
  assign T233 = T18 & T234;
  assign T234 = T168[4'he:4'he];
  assign T282 = reset ? 55'h0 : T235;
  assign T235 = T236 ? io_writeData : regFile_15;
  assign T236 = T18 & T237;
  assign T237 = T168[4'hf:4'hf];
  assign T238 = T174[1'h0:1'h0];
  assign T239 = T174[1'h1:1'h1];
  assign T240 = T174[2'h2:2'h2];
  assign T241 = T174[2'h3:2'h3];
  assign io_full = T242;
  assign T242 = T243 == 16'hffff;
  assign T243 = T3;

  always @(posedge clk) begin
    regRVPipelineRegs_0 <= io_wePipelineReg_0;
    regRVPipelineRegs_1 <= io_wePipelineReg_1;
    regRVPipelineRegs_2 <= io_wePipelineReg_2;
    if(reset) begin
      regPipelineRegs_0 <= 55'h0;
    end else begin
      regPipelineRegs_0 <= io_writePipelineReg_0;
    end
    if(reset) begin
      regPipelineRegs_1 <= 55'h0;
    end else begin
      regPipelineRegs_1 <= io_writePipelineReg_1;
    end
    if(reset) begin
      regPipelineRegs_2 <= 55'h0;
    end else begin
      regPipelineRegs_2 <= io_writePipelineReg_2;
    end
    if(reset) begin
      regFileValid_0 <= 1'h0;
    end else if(T141) begin
      regFileValid_0 <= 1'h0;
    end else if(T9) begin
      regFileValid_0 <= 1'h1;
    end
    if(reset) begin
      writePointer <= 4'h0;
    end else if(T16) begin
      writePointer <= 4'h0;
    end else if(T18) begin
      writePointer <= T15;
    end
    if(reset) begin
      regFileValid_2 <= 1'h0;
    end else if(T30) begin
      regFileValid_2 <= 1'h0;
    end else if(T28) begin
      regFileValid_2 <= 1'h1;
    end
    if(reset) begin
      readPointer <= 4'h0;
    end else if(T37) begin
      readPointer <= 4'h0;
    end else if(io_readIncrement) begin
      readPointer <= T36;
    end
    if(reset) begin
      regFileValid_3 <= 1'h0;
    end else if(T43) begin
      regFileValid_3 <= 1'h0;
    end else if(T41) begin
      regFileValid_3 <= 1'h1;
    end
    if(reset) begin
      regFileValid_4 <= 1'h0;
    end else if(T53) begin
      regFileValid_4 <= 1'h0;
    end else if(T51) begin
      regFileValid_4 <= 1'h1;
    end
    if(reset) begin
      regFileValid_5 <= 1'h0;
    end else if(T59) begin
      regFileValid_5 <= 1'h0;
    end else if(T57) begin
      regFileValid_5 <= 1'h1;
    end
    if(reset) begin
      regFileValid_6 <= 1'h0;
    end else if(T67) begin
      regFileValid_6 <= 1'h0;
    end else if(T65) begin
      regFileValid_6 <= 1'h1;
    end
    if(reset) begin
      regFileValid_7 <= 1'h0;
    end else if(T73) begin
      regFileValid_7 <= 1'h0;
    end else if(T71) begin
      regFileValid_7 <= 1'h1;
    end
    if(reset) begin
      regFileValid_8 <= 1'h0;
    end else if(T85) begin
      regFileValid_8 <= 1'h0;
    end else if(T83) begin
      regFileValid_8 <= 1'h1;
    end
    if(reset) begin
      regFileValid_9 <= 1'h0;
    end else if(T91) begin
      regFileValid_9 <= 1'h0;
    end else if(T89) begin
      regFileValid_9 <= 1'h1;
    end
    if(reset) begin
      regFileValid_10 <= 1'h0;
    end else if(T99) begin
      regFileValid_10 <= 1'h0;
    end else if(T97) begin
      regFileValid_10 <= 1'h1;
    end
    if(reset) begin
      regFileValid_11 <= 1'h0;
    end else if(T105) begin
      regFileValid_11 <= 1'h0;
    end else if(T103) begin
      regFileValid_11 <= 1'h1;
    end
    if(reset) begin
      regFileValid_12 <= 1'h0;
    end else if(T115) begin
      regFileValid_12 <= 1'h0;
    end else if(T113) begin
      regFileValid_12 <= 1'h1;
    end
    if(reset) begin
      regFileValid_13 <= 1'h0;
    end else if(T121) begin
      regFileValid_13 <= 1'h0;
    end else if(T119) begin
      regFileValid_13 <= 1'h1;
    end
    if(reset) begin
      regFileValid_14 <= 1'h0;
    end else if(T129) begin
      regFileValid_14 <= 1'h0;
    end else if(T127) begin
      regFileValid_14 <= 1'h1;
    end
    if(reset) begin
      regFileValid_15 <= 1'h0;
    end else if(T135) begin
      regFileValid_15 <= 1'h0;
    end else if(T133) begin
      regFileValid_15 <= 1'h1;
    end
    if(reset) begin
      regFileValid_1 <= 1'h0;
    end else if(T147) begin
      regFileValid_1 <= 1'h0;
    end else if(T145) begin
      regFileValid_1 <= 1'h1;
    end
    if(reset) begin
      regFile_0 <= 55'h0;
    end else if(T166) begin
      regFile_0 <= io_writeData;
    end
    if(reset) begin
      regFile_1 <= 55'h0;
    end else if(T171) begin
      regFile_1 <= io_writeData;
    end
    if(reset) begin
      regFile_2 <= 55'h0;
    end else if(T177) begin
      regFile_2 <= io_writeData;
    end
    if(reset) begin
      regFile_3 <= 55'h0;
    end else if(T180) begin
      regFile_3 <= io_writeData;
    end
    if(reset) begin
      regFile_4 <= 55'h0;
    end else if(T187) begin
      regFile_4 <= io_writeData;
    end
    if(reset) begin
      regFile_5 <= 55'h0;
    end else if(T190) begin
      regFile_5 <= io_writeData;
    end
    if(reset) begin
      regFile_6 <= 55'h0;
    end else if(T195) begin
      regFile_6 <= io_writeData;
    end
    if(reset) begin
      regFile_7 <= 55'h0;
    end else if(T198) begin
      regFile_7 <= io_writeData;
    end
    if(reset) begin
      regFile_8 <= 55'h0;
    end else if(T207) begin
      regFile_8 <= io_writeData;
    end
    if(reset) begin
      regFile_9 <= 55'h0;
    end else if(T210) begin
      regFile_9 <= io_writeData;
    end
    if(reset) begin
      regFile_10 <= 55'h0;
    end else if(T215) begin
      regFile_10 <= io_writeData;
    end
    if(reset) begin
      regFile_11 <= 55'h0;
    end else if(T218) begin
      regFile_11 <= io_writeData;
    end
    if(reset) begin
      regFile_12 <= 55'h0;
    end else if(T225) begin
      regFile_12 <= io_writeData;
    end
    if(reset) begin
      regFile_13 <= 55'h0;
    end else if(T228) begin
      regFile_13 <= io_writeData;
    end
    if(reset) begin
      regFile_14 <= 55'h0;
    end else if(T233) begin
      regFile_14 <= io_writeData;
    end
    if(reset) begin
      regFile_15 <= 55'h0;
    end else if(T236) begin
      regFile_15 <= io_writeData;
    end
  end
endmodule

module Queue_0(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [54:0] io_enq_bits_x,
    input  io_deq_ready,
    output io_deq_valid,
    output[54:0] io_deq_bits_x,
    output[4:0] io_count
);

  wire[4:0] T0;
  wire[3:0] ptr_diff;
  reg [3:0] R1;
  wire[3:0] T16;
  wire[3:0] T2;
  wire[3:0] T3;
  wire do_deq;
  reg [3:0] R4;
  wire[3:0] T17;
  wire[3:0] T5;
  wire[3:0] T6;
  wire do_enq;
  wire T7;
  wire ptr_match;
  reg  maybe_full;
  wire T18;
  wire T8;
  wire T9;
  wire[54:0] T10;
  wire[54:0] T11;
  reg [54:0] ram [15:0];
  wire[54:0] T12;
  wire T13;
  wire empty;
  wire T14;
  wire T15;
  wire full;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    R1 = {1{1'b0}};
    R4 = {1{1'b0}};
    maybe_full = {1{1'b0}};
    for (initvar = 0; initvar < 16; initvar = initvar+1)
      ram[initvar] = {2{1'b0}};
  end
// synthesis translate_on
`endif

  assign io_count = T0;
  assign T0 = {T7, ptr_diff};
  assign ptr_diff = R4 - R1;
  assign T16 = reset ? 4'h0 : T2;
  assign T2 = do_deq ? T3 : R1;
  assign T3 = R1 + 4'h1;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign T17 = reset ? 4'h0 : T5;
  assign T5 = do_enq ? T6 : R4;
  assign T6 = R4 + 4'h1;
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T7 = maybe_full & ptr_match;
  assign ptr_match = R4 == R1;
  assign T18 = reset ? 1'h0 : T8;
  assign T8 = T9 ? do_enq : maybe_full;
  assign T9 = do_enq != do_deq;
  assign io_deq_bits_x = T10;
  assign T10 = T11[6'h36:1'h0];
  assign T11 = ram[R1];
  assign io_deq_valid = T13;
  assign T13 = empty ^ 1'h1;
  assign empty = ptr_match & T14;
  assign T14 = maybe_full ^ 1'h1;
  assign io_enq_ready = T15;
  assign T15 = full ^ 1'h1;
  assign full = ptr_match & maybe_full;

  always @(posedge clk) begin
    if(reset) begin
      R1 <= 4'h0;
    end else if(do_deq) begin
      R1 <= T3;
    end
    if(reset) begin
      R4 <= 4'h0;
    end else if(do_enq) begin
      R4 <= T6;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T9) begin
      maybe_full <= do_enq;
    end
    if (do_enq)
      ram[R4] <= io_enq_bits_x;
  end
endmodule

module RouterBuffer(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [54:0] io_enq_bits_x,
    input  io_deq_ready,
    output io_deq_valid,
    output[54:0] io_deq_bits_x
);

  wire queue_io_enq_ready;
  wire queue_io_deq_valid;
  wire[54:0] queue_io_deq_bits_x;


  assign io_deq_bits_x = queue_io_deq_bits_x;
  assign io_deq_valid = queue_io_deq_valid;
  assign io_enq_ready = queue_io_enq_ready;
  Queue_0 queue(.clk(clk), .reset(reset),
       .io_enq_ready( queue_io_enq_ready ),
       .io_enq_valid( io_enq_valid ),
       .io_enq_bits_x( io_enq_bits_x ),
       .io_deq_ready( io_deq_ready ),
       .io_deq_valid( queue_io_deq_valid ),
       .io_deq_bits_x( queue_io_deq_bits_x )
       //.io_count(  )
  );
endmodule

module CMeshDOR_0(
    input [15:0] io_inHeadFlit_packetID,
    input  io_inHeadFlit_isTail,
    input  io_inHeadFlit_vcPort,
    input [3:0] io_inHeadFlit_packetType,
    input [1:0] io_inHeadFlit_destination_2,
    input [1:0] io_inHeadFlit_destination_1,
    input [1:0] io_inHeadFlit_destination_0,
    input [2:0] io_inHeadFlit_priorityLevel,
    output[15:0] io_outHeadFlit_packetID,
    output io_outHeadFlit_isTail,
    output io_outHeadFlit_vcPort,
    output[3:0] io_outHeadFlit_packetType,
    output[1:0] io_outHeadFlit_destination_2,
    output[1:0] io_outHeadFlit_destination_1,
    output[1:0] io_outHeadFlit_destination_0,
    output[2:0] io_outHeadFlit_priorityLevel,
    output[2:0] io_result,
    output[1:0] io_vcsAvailable_4,
    output[1:0] io_vcsAvailable_3,
    output[1:0] io_vcsAvailable_2,
    output[1:0] io_vcsAvailable_1,
    output[1:0] io_vcsAvailable_0
);

  wire[1:0] T0;
  wire[1:0] T26;
  wire T1;
  wire[1:0] T2;
  wire[1:0] T27;
  wire T3;
  wire[1:0] T4;
  wire[1:0] T28;
  wire T5;
  wire[1:0] T6;
  wire[1:0] T29;
  wire T7;
  wire[1:0] T8;
  wire[1:0] T30;
  wire T9;
  wire[2:0] T10;
  wire[2:0] resultReduction;
  wire[2:0] T11;
  wire[2:0] dimResults_1;
  wire[2:0] T12;
  wire[2:0] T31;
  wire[1:0] T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire[2:0] dimResults_0;
  wire[2:0] T32;
  wire[1:0] T18;
  wire[1:0] T33;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire[2:0] T34;
  wire T25;


  assign io_vcsAvailable_0 = T0;
  assign T0 = 2'h0 - T26;
  assign T26 = {1'h0, T1};
  assign T1 = io_result == 3'h0;
  assign io_vcsAvailable_1 = T2;
  assign T2 = 2'h0 - T27;
  assign T27 = {1'h0, T3};
  assign T3 = io_result == 3'h1;
  assign io_vcsAvailable_2 = T4;
  assign T4 = 2'h0 - T28;
  assign T28 = {1'h0, T5};
  assign T5 = io_result == 3'h2;
  assign io_vcsAvailable_3 = T6;
  assign T6 = 2'h0 - T29;
  assign T29 = {1'h0, T7};
  assign T7 = io_result == 3'h3;
  assign io_vcsAvailable_4 = T8;
  assign T8 = 2'h0 - T30;
  assign T30 = {1'h0, T9};
  assign T9 = io_result == 3'h4;
  assign io_result = T10;
  assign T10 = T25 ? T34 : resultReduction;
  assign resultReduction = T11;
  assign T11 = T24 ? dimResults_0 : dimResults_1;
  assign dimResults_1 = T12;
  assign T12 = T15 ? 3'h4 : T31;
  assign T31 = {1'h0, T13};
  assign T13 = T14 ? 2'h3 : 2'h0;
  assign T14 = 2'h0 < io_inHeadFlit_destination_1;
  assign T15 = T17 & T16;
  assign T16 = io_inHeadFlit_destination_1 < 2'h0;
  assign T17 = T14 ^ 1'h1;
  assign dimResults_0 = T32;
  assign T32 = {1'h0, T18};
  assign T18 = T21 ? 2'h2 : T33;
  assign T33 = {1'h0, T19};
  assign T19 = T20 ? 1'h1 : 1'h0;
  assign T20 = 2'h0 < io_inHeadFlit_destination_0;
  assign T21 = T23 & T22;
  assign T22 = io_inHeadFlit_destination_0 < 2'h0;
  assign T23 = T20 ^ 1'h1;
  assign T24 = dimResults_0 != 3'h0;
  assign T34 = {1'h0, io_inHeadFlit_destination_2};
  assign T25 = resultReduction == 3'h0;
  assign io_outHeadFlit_priorityLevel = io_inHeadFlit_priorityLevel;
  assign io_outHeadFlit_destination_0 = io_inHeadFlit_destination_0;
  assign io_outHeadFlit_destination_1 = io_inHeadFlit_destination_1;
  assign io_outHeadFlit_destination_2 = io_inHeadFlit_destination_2;
  assign io_outHeadFlit_packetType = io_inHeadFlit_packetType;
  assign io_outHeadFlit_vcPort = io_inHeadFlit_vcPort;
  assign io_outHeadFlit_isTail = io_inHeadFlit_isTail;
  assign io_outHeadFlit_packetID = io_inHeadFlit_packetID;
endmodule

module VCRouterStateManagement(input clk, input reset,
    input  io_inputBufferValid,
    input  io_routingComplete,
    input  io_inputBufferIsTail,
    input  io_vcAllocGranted,
    input  io_swAllocGranted,
    input  io_creditsAvail,
    input  io_outputReady,
    output[2:0] io_currentState
);

  reg [2:0] curState;
  wire[2:0] T56;
  wire[2:0] T0;
  wire[2:0] T1;
  wire[2:0] T2;
  wire[2:0] T3;
  wire[2:0] T4;
  wire[2:0] T5;
  wire[2:0] T6;
  wire[2:0] T7;
  wire[2:0] T8;
  wire[2:0] T9;
  wire[2:0] T10;
  wire[2:0] T11;
  wire[2:0] T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    curState = {1{1'b0}};
  end
// synthesis translate_on
`endif

  assign io_currentState = curState;
  assign T56 = reset ? 3'h0 : T0;
  assign T0 = T54 ? 3'h5 : T1;
  assign T1 = T49 ? 3'h4 : T2;
  assign T2 = T46 ? 3'h5 : T3;
  assign T3 = T43 ? 3'h4 : T4;
  assign T4 = T37 ? 3'h0 : T5;
  assign T5 = T35 ? 3'h3 : T6;
  assign T6 = T30 ? 3'h4 : T7;
  assign T7 = T28 ? 3'h2 : T8;
  assign T8 = T23 ? 3'h3 : T9;
  assign T9 = T21 ? 3'h1 : T10;
  assign T10 = T17 ? 3'h2 : T11;
  assign T11 = T15 ? 3'h0 : T12;
  assign T12 = T13 ? 3'h1 : curState;
  assign T13 = T14 & io_inputBufferValid;
  assign T14 = curState == 3'h0;
  assign T15 = T14 & T16;
  assign T16 = io_inputBufferValid ^ 1'h1;
  assign T17 = T18 & io_routingComplete;
  assign T18 = T20 & T19;
  assign T19 = curState == 3'h1;
  assign T20 = T14 ^ 1'h1;
  assign T21 = T18 & T22;
  assign T22 = io_routingComplete ^ 1'h1;
  assign T23 = T24 & io_vcAllocGranted;
  assign T24 = T26 & T25;
  assign T25 = curState == 3'h2;
  assign T26 = T27 ^ 1'h1;
  assign T27 = T14 | T19;
  assign T28 = T24 & T29;
  assign T29 = io_vcAllocGranted ^ 1'h1;
  assign T30 = T31 & io_swAllocGranted;
  assign T31 = T33 & T32;
  assign T32 = curState == 3'h3;
  assign T33 = T34 ^ 1'h1;
  assign T34 = T27 | T25;
  assign T35 = T31 & T36;
  assign T36 = io_swAllocGranted ^ 1'h1;
  assign T37 = T39 & T38;
  assign T38 = io_inputBufferIsTail & io_creditsAvail;
  assign T39 = T41 & T40;
  assign T40 = curState == 3'h4;
  assign T41 = T42 ^ 1'h1;
  assign T42 = T34 | T32;
  assign T43 = T39 & T44;
  assign T44 = T45 & io_creditsAvail;
  assign T45 = T38 ^ 1'h1;
  assign T46 = T39 & T47;
  assign T47 = T48 ^ 1'h1;
  assign T48 = T38 | io_creditsAvail;
  assign T49 = T50 & io_creditsAvail;
  assign T50 = T52 & T51;
  assign T51 = curState == 3'h5;
  assign T52 = T53 ^ 1'h1;
  assign T53 = T42 | T40;
  assign T54 = T50 & T55;
  assign T55 = io_creditsAvail ^ 1'h1;

  always @(posedge clk) begin
    if(reset) begin
      curState <= 3'h0;
    end else if(T54) begin
      curState <= 3'h5;
    end else if(T49) begin
      curState <= 3'h4;
    end else if(T46) begin
      curState <= 3'h5;
    end else if(T43) begin
      curState <= 3'h4;
    end else if(T37) begin
      curState <= 3'h0;
    end else if(T35) begin
      curState <= 3'h3;
    end else if(T30) begin
      curState <= 3'h4;
    end else if(T28) begin
      curState <= 3'h2;
    end else if(T23) begin
      curState <= 3'h3;
    end else if(T21) begin
      curState <= 3'h1;
    end else if(T17) begin
      curState <= 3'h2;
    end else if(T15) begin
      curState <= 3'h0;
    end else if(T13) begin
      curState <= 3'h1;
    end
  end
endmodule

module MuxN_0(
    input [54:0] io_ins_1_x,
    input [54:0] io_ins_0_x,
    input  io_sel,
    output[54:0] io_out_x
);

  wire[54:0] T0;
  wire T1;


  assign io_out_x = T0;
  assign T0 = T1 ? io_ins_1_x : io_ins_0_x;
  assign T1 = io_sel;
endmodule

module ReplaceVCPort(
    input [54:0] io_oldFlit_x,
    input  io_newVCPort,
    output[54:0] io_newFlit_x
);

  wire T0;
  wire T1;
  wire[54:0] T2;
  wire[54:0] T3;
  wire[53:0] T4;
  wire[53:0] T5;
  wire[36:0] T6;
  wire[35:0] T7;
  wire[31:0] b_payload;
  wire[31:0] T8;
  wire[53:0] T9;
  wire[3:0] b_flitID;
  wire[3:0] T10;
  wire[53:0] T11;
  wire b_vcPort;
  wire[16:0] T12;
  wire b_isTail;
  wire T13;
  wire[53:0] T14;
  wire[15:0] b_packetID;
  wire[15:0] T15;
  wire[53:0] T16;
  wire[54:0] T17;
  wire[54:0] T18;
  wire[31:0] T19;
  wire[30:0] T20;
  wire[30:0] T21;
  wire[8:0] T22;
  wire[4:0] T23;
  wire[2:0] h_priorityLevel;
  wire[1:0] h_destination_0;
  wire[1:0] T24;
  wire[30:0] T25;
  wire[3:0] T26;
  wire[1:0] h_destination_1;
  wire[1:0] T27;
  wire[30:0] T28;
  wire[1:0] h_destination_2;
  wire[1:0] T29;
  wire[30:0] T30;
  wire[21:0] T31;
  wire[4:0] T32;
  wire[3:0] h_packetType;
  wire[3:0] T33;
  wire[30:0] T34;
  wire h_vcPort;
  wire[16:0] T35;
  wire h_isTail;
  wire T36;
  wire[30:0] T37;
  wire[15:0] h_packetID;
  wire[15:0] T38;
  wire[30:0] T39;
  wire[54:0] flitVCMux_io_out_x;


`ifndef SYNTHESIS
// synthesis translate_off
  assign h_priorityLevel = {1{1'b0}};
// synthesis translate_on
`endif
  assign T0 = T1 == 1'h1;
  assign T1 = io_oldFlit_x[1'h0:1'h0];
  assign T2 = T3;
  assign T3 = {T4, 1'h0};
  assign T4 = T5;
  assign T5 = {T12, T6};
  assign T6 = {b_vcPort, T7};
  assign T7 = {b_flitID, b_payload};
  assign b_payload = T8;
  assign T8 = T9[5'h1f:1'h0];
  assign T9 = io_oldFlit_x[6'h36:1'h1];
  assign b_flitID = T10;
  assign T10 = T11[6'h23:6'h20];
  assign T11 = io_oldFlit_x[6'h36:1'h1];
  assign b_vcPort = io_newVCPort;
  assign T12 = {b_packetID, b_isTail};
  assign b_isTail = T13;
  assign T13 = T14[6'h25:6'h25];
  assign T14 = io_oldFlit_x[6'h36:1'h1];
  assign b_packetID = T15;
  assign T15 = T16[6'h35:6'h26];
  assign T16 = io_oldFlit_x[6'h36:1'h1];
  assign T17 = T18;
  assign T18 = {23'h0, T19};
  assign T19 = {T20, 1'h1};
  assign T20 = T21;
  assign T21 = {T31, T22};
  assign T22 = {T26, T23};
  assign T23 = {h_destination_0, h_priorityLevel};
  assign h_destination_0 = T24;
  assign T24 = T25[3'h4:2'h3];
  assign T25 = io_oldFlit_x[5'h1f:1'h1];
  assign T26 = {h_destination_2, h_destination_1};
  assign h_destination_1 = T27;
  assign T27 = T28[3'h6:3'h5];
  assign T28 = io_oldFlit_x[5'h1f:1'h1];
  assign h_destination_2 = T29;
  assign T29 = T30[4'h8:3'h7];
  assign T30 = io_oldFlit_x[5'h1f:1'h1];
  assign T31 = {T35, T32};
  assign T32 = {h_vcPort, h_packetType};
  assign h_packetType = T33;
  assign T33 = T34[4'hc:4'h9];
  assign T34 = io_oldFlit_x[5'h1f:1'h1];
  assign h_vcPort = io_newVCPort;
  assign T35 = {h_packetID, h_isTail};
  assign h_isTail = T36;
  assign T36 = T37[4'he:4'he];
  assign T37 = io_oldFlit_x[5'h1f:1'h1];
  assign h_packetID = T38;
  assign T38 = T39[5'h1e:4'hf];
  assign T39 = io_oldFlit_x[5'h1f:1'h1];
  assign io_newFlit_x = flitVCMux_io_out_x;
  MuxN_0 flitVCMux(
       .io_ins_1_x( T17 ),
       .io_ins_0_x( T2 ),
       .io_sel( T0 ),
       .io_out_x( flitVCMux_io_out_x )
  );
endmodule

module Flit2FlitBundle(
    input [54:0] io_inFlit_x,
    output[15:0] io_outHead_packetID,
    output io_outHead_isTail,
    output io_outHead_vcPort,
    output[3:0] io_outHead_packetType,
    output[1:0] io_outHead_destination_2,
    output[1:0] io_outHead_destination_1,
    output[1:0] io_outHead_destination_0,
    output[2:0] io_outHead_priorityLevel,
    output[15:0] io_outBody_packetID,
    output io_outBody_isTail,
    output io_outBody_vcPort,
    output[3:0] io_outBody_flitID,
    output[31:0] io_outBody_payload
);

  wire[31:0] T0;
  wire[53:0] T1;
  wire[3:0] T2;
  wire T3;
  wire T4;
  wire[15:0] T5;
  wire[2:0] T6;
  wire[30:0] T7;
  wire[1:0] T8;
  wire[1:0] T9;
  wire[1:0] T10;
  wire[3:0] T11;
  wire T12;
  wire T13;
  wire[15:0] T14;


  assign io_outBody_payload = T0;
  assign T0 = T1[5'h1f:1'h0];
  assign T1 = io_inFlit_x[6'h36:1'h1];
  assign io_outBody_flitID = T2;
  assign T2 = T1[6'h23:6'h20];
  assign io_outBody_vcPort = T3;
  assign T3 = T1[6'h24:6'h24];
  assign io_outBody_isTail = T4;
  assign T4 = T1[6'h25:6'h25];
  assign io_outBody_packetID = T5;
  assign T5 = T1[6'h35:6'h26];
  assign io_outHead_priorityLevel = T6;
  assign T6 = T7[2'h2:1'h0];
  assign T7 = io_inFlit_x[5'h1f:1'h1];
  assign io_outHead_destination_0 = T8;
  assign T8 = T7[3'h4:2'h3];
  assign io_outHead_destination_1 = T9;
  assign T9 = T7[3'h6:3'h5];
  assign io_outHead_destination_2 = T10;
  assign T10 = T7[4'h8:3'h7];
  assign io_outHead_packetType = T11;
  assign T11 = T7[4'hc:4'h9];
  assign io_outHead_vcPort = T12;
  assign T12 = T7[4'hd:4'hd];
  assign io_outHead_isTail = T13;
  assign T13 = T7[4'he:4'he];
  assign io_outHead_packetID = T14;
  assign T14 = T7[5'h1e:4'hf];
endmodule

module CreditCon(input clk, input reset,
    input  io_inCredit_grant,
    input  io_inConsume,
    output io_outCredit,
    output io_almostOut
);

  reg[0:0] T0;
  wire T1;
  wire T2;
  reg [4:0] credCount;
  wire[4:0] T22;
  wire[4:0] T3;
  wire[4:0] T4;
  wire[4:0] T5;
  wire[4:0] T6;
  wire[4:0] T23;
  wire T7;
  wire T8;
  wire[4:0] T9;
  wire[4:0] T24;
  wire T10;
  wire[4:0] T11;
  wire[4:0] T25;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire[4:0] T16;
  wire[4:0] T26;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    T0 = 1'b0;
    credCount = {1{1'b0}};
  end
// synthesis translate_on
`endif

  assign T1 = T2 | reset;
  assign T2 = credCount <= 5'h10;
  assign T22 = reset ? 5'h10 : T3;
  assign T3 = T18 ? T16 : T4;
  assign T4 = T13 ? T9 : T5;
  assign T5 = T8 ? T6 : credCount;
  assign T6 = credCount - T23;
  assign T23 = {4'h0, T7};
  assign T7 = io_inConsume;
  assign T8 = credCount == 5'h10;
  assign T9 = T11 - T24;
  assign T24 = {4'h0, T10};
  assign T10 = io_inConsume;
  assign T11 = credCount + T25;
  assign T25 = {4'h0, T12};
  assign T12 = io_inCredit_grant;
  assign T13 = T15 & T14;
  assign T14 = 5'h1 < credCount;
  assign T15 = T8 ^ 1'h1;
  assign T16 = credCount + T26;
  assign T26 = {4'h0, T17};
  assign T17 = io_inCredit_grant;
  assign T18 = T19 ^ 1'h1;
  assign T19 = T8 | T14;
  assign io_almostOut = T20;
  assign T20 = credCount == 5'h2;
  assign io_outCredit = T21;
  assign T21 = 5'h1 < credCount;

  always @(posedge clk) begin
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T0 <= 1'b1;
  if(!T1 && T0 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "CreditCon: Exceeded max credits");
    $finish;
  end
// synthesis translate_on
`endif
    if(reset) begin
      credCount <= 5'h10;
    end else if(T18) begin
      credCount <= T16;
    end else if(T13) begin
      credCount <= T9;
    end else if(T8) begin
      credCount <= T6;
    end
  end
endmodule

module MuxN_1(
    input  io_ins_1,
    input  io_ins_0,
    input  io_sel,
    output io_out
);

  wire T0;
  wire T1;


  assign io_out = T0;
  assign T0 = T1 ? io_ins_1 : io_ins_0;
  assign T1 = io_sel;
endmodule

module SimpleVCRouter_0((* gated_clock = "true" *) input clk, input reset,
    input [54:0] io_inChannels_4_flit_x,
    input  io_inChannels_4_flitValid,
    output io_inChannels_4_credit_1_grant,
    output io_inChannels_4_credit_0_grant,
    input [54:0] io_inChannels_3_flit_x,
    input  io_inChannels_3_flitValid,
    output io_inChannels_3_credit_1_grant,
    output io_inChannels_3_credit_0_grant,
    input [54:0] io_inChannels_2_flit_x,
    input  io_inChannels_2_flitValid,
    output io_inChannels_2_credit_1_grant,
    output io_inChannels_2_credit_0_grant,
    input [54:0] io_inChannels_1_flit_x,
    input  io_inChannels_1_flitValid,
    output io_inChannels_1_credit_1_grant,
    output io_inChannels_1_credit_0_grant,
    input [54:0] io_inChannels_0_flit_x,
    input  io_inChannels_0_flitValid,
    output io_inChannels_0_credit_1_grant,
    output io_inChannels_0_credit_0_grant,
    output[54:0] io_outChannels_4_flit_x,
    output io_outChannels_4_flitValid,
    input  io_outChannels_4_credit_1_grant,
    input  io_outChannels_4_credit_0_grant,
    output[54:0] io_outChannels_3_flit_x,
    output io_outChannels_3_flitValid,
    input  io_outChannels_3_credit_1_grant,
    input  io_outChannels_3_credit_0_grant,
    output[54:0] io_outChannels_2_flit_x,
    output io_outChannels_2_flitValid,
    input  io_outChannels_2_credit_1_grant,
    input  io_outChannels_2_credit_0_grant,
    output[54:0] io_outChannels_1_flit_x,
    output io_outChannels_1_flitValid,
    input  io_outChannels_1_credit_1_grant,
    input  io_outChannels_1_credit_0_grant,
    output[54:0] io_outChannels_0_flit_x,
    output io_outChannels_0_flitValid,
    input  io_outChannels_0_credit_1_grant,
    input  io_outChannels_0_credit_0_grant,
    //output[31:0] io_counters_1_counterVal
    //output[7:0] io_counters_1_counterIndex
    output[31:0] io_counters_0_counterVal
    //output[7:0] io_counters_0_counterIndex
    //input  io_bypass
);

  reg[0:0] T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  wire[53:0] T8;
  wire T9;
  wire[30:0] T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  reg[0:0] T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  reg[0:0] T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire[53:0] T30;
  wire T31;
  wire[30:0] T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  reg[0:0] T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  reg[0:0] T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire[53:0] T52;
  wire T53;
  wire[30:0] T54;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  reg[0:0] T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  reg[0:0] T66;
  wire T67;
  wire T68;
  wire T69;
  wire T70;
  wire T71;
  wire T72;
  wire T73;
  wire[53:0] T74;
  wire T75;
  wire[30:0] T76;
  wire T77;
  wire T78;
  wire T79;
  wire T80;
  wire T81;
  wire T82;
  reg[0:0] T83;
  wire T84;
  wire T85;
  wire T86;
  wire T87;
  reg[0:0] T88;
  wire T89;
  wire T90;
  wire T91;
  wire T92;
  wire T93;
  wire T94;
  wire T95;
  wire[53:0] T96;
  wire T97;
  wire[30:0] T98;
  wire T99;
  wire T100;
  wire T101;
  wire T102;
  wire T103;
  wire T104;
  reg[0:0] T105;
  wire T106;
  wire T107;
  wire T108;
  wire T109;
  reg[0:0] T110;
  wire T111;
  wire T112;
  wire T113;
  wire T114;
  wire T115;
  wire T116;
  wire T117;
  wire[53:0] T118;
  wire T119;
  wire[30:0] T120;
  wire T121;
  wire T122;
  wire T123;
  wire T124;
  wire T125;
  wire T126;
  reg[0:0] T127;
  wire T128;
  wire T129;
  wire T130;
  wire T131;
  reg[0:0] T132;
  wire T133;
  wire T134;
  wire T135;
  wire T136;
  wire T137;
  wire T138;
  wire T139;
  wire[53:0] T140;
  wire T141;
  wire[30:0] T142;
  wire T143;
  wire T144;
  wire T145;
  wire T146;
  wire T147;
  wire T148;
  reg[0:0] T149;
  wire T150;
  wire T151;
  wire T152;
  wire T153;
  reg[0:0] T154;
  wire T155;
  wire T156;
  wire T157;
  wire T158;
  wire T159;
  wire T160;
  wire T161;
  wire[53:0] T162;
  wire T163;
  wire[30:0] T164;
  wire T165;
  wire T166;
  wire T167;
  wire T168;
  wire T169;
  wire T170;
  reg[0:0] T171;
  wire T172;
  wire T173;
  wire T174;
  wire T175;
  reg[0:0] T176;
  wire T177;
  wire T178;
  wire T179;
  wire T180;
  wire T181;
  wire T182;
  wire T183;
  wire[53:0] T184;
  wire T185;
  wire[30:0] T186;
  wire T187;
  wire T188;
  wire T189;
  wire T190;
  wire T191;
  wire T192;
  reg[0:0] T193;
  wire T194;
  wire T195;
  wire T196;
  wire T197;
  reg[0:0] T198;
  wire T199;
  wire T200;
  wire T201;
  wire T202;
  wire T203;
  wire T204;
  wire T205;
  wire[53:0] T206;
  wire T207;
  wire[30:0] T208;
  wire T209;
  wire T210;
  wire T211;
  wire T212;
  wire T213;
  wire T214;
  reg[0:0] T215;
  wire T216;
  wire T217;
  wire T218;
  wire T219;
  wire T220;
  wire T221;
  wire T222;
  wire T223;
  wire T224;
  wire[53:0] T225;
  wire T226;
  wire[30:0] T227;
  wire T228;
  wire T229;
  wire T230;
  wire T231;
  wire T232;
  wire T233;
  wire T234;
  wire T235;
  wire T236;
  wire[53:0] T237;
  wire T238;
  wire[30:0] T239;
  wire T240;
  wire T241;
  wire T242;
  wire T243;
  wire T244;
  wire T245;
  wire T246;
  wire T247;
  wire T248;
  wire[53:0] T249;
  wire T250;
  wire[30:0] T251;
  wire T252;
  wire T253;
  wire T254;
  wire T255;
  wire T256;
  wire T257;
  wire T258;
  wire T259;
  wire T260;
  wire[53:0] T261;
  wire T262;
  wire[30:0] T263;
  wire T264;
  wire T265;
  wire T266;
  wire T267;
  wire T268;
  wire T269;
  wire T270;
  wire T271;
  wire T272;
  wire[53:0] T273;
  wire T274;
  wire[30:0] T275;
  wire T276;
  wire T277;
  wire T278;
  wire T279;
  wire[54:0] T280;
  wire[54:0] T281;
  wire T3112;
  reg [54:0] R282;
  wire[54:0] T3113;
  wire[54:0] T283;
  wire[54:0] T3114;
  wire T284;
  wire T285;
  wire[54:0] T286;
  wire[54:0] T287;
  wire T288;
  wire T289;
  wire[1:0] T290;
  wire[1:0] T291;
  wire[1:0] T292;
  wire T293;
  wire[2:0] T294;
  reg [2:0] R295;
  wire[2:0] T3115;
  wire[1:0] T296;
  wire T297;
  wire T298;
  wire T299;
  wire T300;
  wire T301;
  wire T302;
  wire T303;
  wire T304;
  wire creditConsReady_0_0;
  wire creditConsReady_1_0;
  wire T305;
  wire[2:0] T306;
  wire T307;
  wire creditConsReady_2_0;
  wire creditConsReady_3_0;
  wire T308;
  wire T309;
  wire creditConsReady_4_0;
  wire T310;
  wire T311;
  wire T312;
  wire T313;
  wire creditConsReady_0_1;
  wire creditConsReady_1_1;
  wire T314;
  wire T315;
  wire creditConsReady_2_1;
  wire creditConsReady_3_1;
  wire T316;
  wire T317;
  wire creditConsReady_4_1;
  wire T318;
  wire T319;
  wire T3116;
  wire T320;
  wire T321;
  wire[3:0] T322;
  wire[3:0] T323;
  wire[3:0] T324;
  wire T325;
  wire[2:0] T326;
  wire[3:0] T327;
  wire T328;
  wire T329;
  wire T330;
  wire T331;
  wire T332;
  wire T333;
  wire T334;
  wire[2:0] T335;
  wire T336;
  wire T337;
  wire T338;
  wire T339;
  wire T340;
  wire T341;
  wire T342;
  wire T343;
  wire[53:0] T344;
  wire T345;
  wire[30:0] T346;
  wire T347;
  wire T348;
  reg  R349;
  wire T3117;
  wire[2:0] T350;
  wire[30:0] T351;
  wire[54:0] T352;
  wire[1:0] T353;
  wire[1:0] T354;
  wire[1:0] T355;
  wire[3:0] T356;
  wire T357;
  wire T358;
  wire[15:0] T359;
  wire T360;
  wire T361;
  wire T362;
  wire T363;
  wire T364;
  wire T365;
  wire T366;
  wire T367;
  wire T368;
  wire T369;
  wire T370;
  wire T371;
  wire T372;
  wire T373;
  wire T374;
  wire T375;
  wire T376;
  wire T377;
  wire T378;
  wire T379;
  wire T380;
  wire T381;
  wire T382;
  wire T383;
  wire T384;
  wire T385;
  wire T386;
  wire T387;
  wire[54:0] T3118;
  wire[30:0] T388;
  wire[30:0] T389;
  wire[8:0] T390;
  wire[4:0] T391;
  wire[3:0] T392;
  wire[21:0] T393;
  wire[4:0] T394;
  wire[16:0] T395;
  wire T396;
  wire T397;
  wire T398;
  wire T399;
  wire flitsAreTail_9;
  wire T400;
  wire T401;
  wire T402;
  wire T403;
  wire[53:0] T404;
  wire T405;
  wire[30:0] T406;
  wire T407;
  wire T408;
  wire T409;
  wire T410;
  wire T411;
  wire[54:0] T412;
  wire[54:0] T413;
  wire T414;
  wire T415;
  wire T416;
  wire T417;
  wire T418;
  wire T419;
  wire T420;
  wire T421;
  wire T422;
  wire T423;
  wire[54:0] T424;
  wire[54:0] T425;
  wire T3119;
  reg [54:0] R426;
  wire[54:0] T3120;
  wire[54:0] T427;
  wire[54:0] T3121;
  wire T428;
  wire T429;
  wire[54:0] T430;
  wire[54:0] T431;
  wire T432;
  wire T433;
  wire[1:0] T434;
  wire[1:0] T435;
  wire[1:0] T436;
  wire T437;
  wire[2:0] T438;
  reg [2:0] R439;
  wire[2:0] T3122;
  wire[1:0] T440;
  wire T441;
  wire T442;
  wire T443;
  wire T444;
  wire T445;
  wire T446;
  wire T447;
  wire T448;
  wire T449;
  wire[2:0] T450;
  wire T451;
  wire T452;
  wire T453;
  wire T454;
  wire T455;
  wire T456;
  wire T457;
  wire T458;
  wire T459;
  wire T460;
  wire T461;
  wire T462;
  wire T463;
  wire T3123;
  wire T464;
  wire T465;
  wire[3:0] T466;
  wire[3:0] T467;
  wire[3:0] T468;
  wire T469;
  wire[2:0] T470;
  wire[3:0] T471;
  wire T472;
  wire T473;
  wire T474;
  wire T475;
  wire T476;
  wire T477;
  wire T478;
  wire[2:0] T479;
  wire T480;
  wire T481;
  wire T482;
  wire T483;
  wire T484;
  wire T485;
  wire T486;
  wire T487;
  wire[53:0] T488;
  wire T489;
  wire[30:0] T490;
  wire T491;
  wire T492;
  reg  R493;
  wire T3124;
  wire[2:0] T494;
  wire[30:0] T495;
  wire[54:0] T496;
  wire[1:0] T497;
  wire[1:0] T498;
  wire[1:0] T499;
  wire[3:0] T500;
  wire T501;
  wire T502;
  wire[15:0] T503;
  wire T504;
  wire T505;
  wire T506;
  wire T507;
  wire T508;
  wire T509;
  wire T510;
  wire T511;
  wire T512;
  wire T513;
  wire T514;
  wire T515;
  wire T516;
  wire T517;
  wire T518;
  wire T519;
  wire T520;
  wire T521;
  wire T522;
  wire T523;
  wire T524;
  wire T525;
  wire T526;
  wire T527;
  wire T528;
  wire T529;
  wire T530;
  wire T531;
  wire[54:0] T3125;
  wire[30:0] T532;
  wire[30:0] T533;
  wire[8:0] T534;
  wire[4:0] T535;
  wire[3:0] T536;
  wire[21:0] T537;
  wire[4:0] T538;
  wire[16:0] T539;
  wire T540;
  wire T541;
  wire T542;
  wire T543;
  wire flitsAreTail_8;
  wire T544;
  wire T545;
  wire T546;
  wire T547;
  wire[53:0] T548;
  wire T549;
  wire[30:0] T550;
  wire T551;
  wire T552;
  wire T553;
  wire T554;
  wire T555;
  wire[54:0] T556;
  wire[54:0] T557;
  wire T558;
  wire T559;
  wire T560;
  wire T561;
  wire T562;
  wire T563;
  wire T564;
  wire T565;
  wire T566;
  wire T567;
  wire[54:0] T568;
  wire[54:0] T569;
  wire T3126;
  reg [54:0] R570;
  wire[54:0] T3127;
  wire[54:0] T571;
  wire[54:0] T3128;
  wire T572;
  wire T573;
  wire[54:0] T574;
  wire[54:0] T575;
  wire T576;
  wire T577;
  wire[1:0] T578;
  wire[1:0] T579;
  wire[1:0] T580;
  wire T581;
  wire[2:0] T582;
  reg [2:0] R583;
  wire[2:0] T3129;
  wire[1:0] T584;
  wire T585;
  wire T586;
  wire T587;
  wire T588;
  wire T589;
  wire T590;
  wire T591;
  wire T592;
  wire T593;
  wire[2:0] T594;
  wire T595;
  wire T596;
  wire T597;
  wire T598;
  wire T599;
  wire T600;
  wire T601;
  wire T602;
  wire T603;
  wire T604;
  wire T605;
  wire T606;
  wire T607;
  wire T3130;
  wire T608;
  wire T609;
  wire[3:0] T610;
  wire[3:0] T611;
  wire[3:0] T612;
  wire T613;
  wire[2:0] T614;
  wire[3:0] T615;
  wire T616;
  wire T617;
  wire T618;
  wire T619;
  wire T620;
  wire T621;
  wire T622;
  wire[2:0] T623;
  wire T624;
  wire T625;
  wire T626;
  wire T627;
  wire T628;
  wire T629;
  wire T630;
  wire T631;
  wire[53:0] T632;
  wire T633;
  wire[30:0] T634;
  wire T635;
  wire T636;
  reg  R637;
  wire T3131;
  wire[2:0] T638;
  wire[30:0] T639;
  wire[54:0] T640;
  wire[1:0] T641;
  wire[1:0] T642;
  wire[1:0] T643;
  wire[3:0] T644;
  wire T645;
  wire T646;
  wire[15:0] T647;
  wire T648;
  wire T649;
  wire T650;
  wire T651;
  wire T652;
  wire T653;
  wire T654;
  wire T655;
  wire T656;
  wire T657;
  wire T658;
  wire T659;
  wire T660;
  wire T661;
  wire T662;
  wire T663;
  wire T664;
  wire T665;
  wire T666;
  wire T667;
  wire T668;
  wire T669;
  wire T670;
  wire T671;
  wire T672;
  wire T673;
  wire T674;
  wire T675;
  wire[54:0] T3132;
  wire[30:0] T676;
  wire[30:0] T677;
  wire[8:0] T678;
  wire[4:0] T679;
  wire[3:0] T680;
  wire[21:0] T681;
  wire[4:0] T682;
  wire[16:0] T683;
  wire T684;
  wire T685;
  wire T686;
  wire T687;
  wire flitsAreTail_7;
  wire T688;
  wire T689;
  wire T690;
  wire T691;
  wire[53:0] T692;
  wire T693;
  wire[30:0] T694;
  wire T695;
  wire T696;
  wire T697;
  wire T698;
  wire T699;
  wire[54:0] T700;
  wire[54:0] T701;
  wire T702;
  wire T703;
  wire T704;
  wire T705;
  wire T706;
  wire T707;
  wire T708;
  wire T709;
  wire T710;
  wire T711;
  wire[54:0] T712;
  wire[54:0] T713;
  wire T3133;
  reg [54:0] R714;
  wire[54:0] T3134;
  wire[54:0] T715;
  wire[54:0] T3135;
  wire T716;
  wire T717;
  wire[54:0] T718;
  wire[54:0] T719;
  wire T720;
  wire T721;
  wire[1:0] T722;
  wire[1:0] T723;
  wire[1:0] T724;
  wire T725;
  wire[2:0] T726;
  reg [2:0] R727;
  wire[2:0] T3136;
  wire[1:0] T728;
  wire T729;
  wire T730;
  wire T731;
  wire T732;
  wire T733;
  wire T734;
  wire T735;
  wire T736;
  wire T737;
  wire[2:0] T738;
  wire T739;
  wire T740;
  wire T741;
  wire T742;
  wire T743;
  wire T744;
  wire T745;
  wire T746;
  wire T747;
  wire T748;
  wire T749;
  wire T750;
  wire T751;
  wire T3137;
  wire T752;
  wire T753;
  wire[3:0] T754;
  wire[3:0] T755;
  wire[3:0] T756;
  wire T757;
  wire[2:0] T758;
  wire[3:0] T759;
  wire T760;
  wire T761;
  wire T762;
  wire T763;
  wire T764;
  wire T765;
  wire T766;
  wire[2:0] T767;
  wire T768;
  wire T769;
  wire T770;
  wire T771;
  wire T772;
  wire T773;
  wire T774;
  wire T775;
  wire[53:0] T776;
  wire T777;
  wire[30:0] T778;
  wire T779;
  wire T780;
  reg  R781;
  wire T3138;
  wire[2:0] T782;
  wire[30:0] T783;
  wire[54:0] T784;
  wire[1:0] T785;
  wire[1:0] T786;
  wire[1:0] T787;
  wire[3:0] T788;
  wire T789;
  wire T790;
  wire[15:0] T791;
  wire T792;
  wire T793;
  wire T794;
  wire T795;
  wire T796;
  wire T797;
  wire T798;
  wire T799;
  wire T800;
  wire T801;
  wire T802;
  wire T803;
  wire T804;
  wire T805;
  wire T806;
  wire T807;
  wire T808;
  wire T809;
  wire T810;
  wire T811;
  wire T812;
  wire T813;
  wire T814;
  wire T815;
  wire T816;
  wire T817;
  wire T818;
  wire T819;
  wire[54:0] T3139;
  wire[30:0] T820;
  wire[30:0] T821;
  wire[8:0] T822;
  wire[4:0] T823;
  wire[3:0] T824;
  wire[21:0] T825;
  wire[4:0] T826;
  wire[16:0] T827;
  wire T828;
  wire T829;
  wire T830;
  wire T831;
  wire flitsAreTail_6;
  wire T832;
  wire T833;
  wire T834;
  wire T835;
  wire[53:0] T836;
  wire T837;
  wire[30:0] T838;
  wire T839;
  wire T840;
  wire T841;
  wire T842;
  wire T843;
  wire[54:0] T844;
  wire[54:0] T845;
  wire T846;
  wire T847;
  wire T848;
  wire T849;
  wire T850;
  wire T851;
  wire T852;
  wire T853;
  wire T854;
  wire T855;
  wire[54:0] T856;
  wire[54:0] T857;
  wire T3140;
  reg [54:0] R858;
  wire[54:0] T3141;
  wire[54:0] T859;
  wire[54:0] T3142;
  wire T860;
  wire T861;
  wire[54:0] T862;
  wire[54:0] T863;
  wire T864;
  wire T865;
  wire[1:0] T866;
  wire[1:0] T867;
  wire[1:0] T868;
  wire T869;
  wire[2:0] T870;
  reg [2:0] R871;
  wire[2:0] T3143;
  wire[1:0] T872;
  wire T873;
  wire T874;
  wire T875;
  wire T876;
  wire T877;
  wire T878;
  wire T879;
  wire T880;
  wire T881;
  wire[2:0] T882;
  wire T883;
  wire T884;
  wire T885;
  wire T886;
  wire T887;
  wire T888;
  wire T889;
  wire T890;
  wire T891;
  wire T892;
  wire T893;
  wire T894;
  wire T895;
  wire T3144;
  wire T896;
  wire T897;
  wire[3:0] T898;
  wire[3:0] T899;
  wire[3:0] T900;
  wire T901;
  wire[2:0] T902;
  wire[3:0] T903;
  wire T904;
  wire T905;
  wire T906;
  wire T907;
  wire T908;
  wire T909;
  wire T910;
  wire[2:0] T911;
  wire T912;
  wire T913;
  wire T914;
  wire T915;
  wire T916;
  wire T917;
  wire T918;
  wire T919;
  wire[53:0] T920;
  wire T921;
  wire[30:0] T922;
  wire T923;
  wire T924;
  reg  R925;
  wire T3145;
  wire[2:0] T926;
  wire[30:0] T927;
  wire[54:0] T928;
  wire[1:0] T929;
  wire[1:0] T930;
  wire[1:0] T931;
  wire[3:0] T932;
  wire T933;
  wire T934;
  wire[15:0] T935;
  wire T936;
  wire T937;
  wire T938;
  wire T939;
  wire T940;
  wire T941;
  wire T942;
  wire T943;
  wire T944;
  wire T945;
  wire T946;
  wire T947;
  wire T948;
  wire T949;
  wire T950;
  wire T951;
  wire T952;
  wire T953;
  wire T954;
  wire T955;
  wire T956;
  wire T957;
  wire T958;
  wire T959;
  wire T960;
  wire T961;
  wire T962;
  wire T963;
  wire[54:0] T3146;
  wire[30:0] T964;
  wire[30:0] T965;
  wire[8:0] T966;
  wire[4:0] T967;
  wire[3:0] T968;
  wire[21:0] T969;
  wire[4:0] T970;
  wire[16:0] T971;
  wire T972;
  wire T973;
  wire T974;
  wire T975;
  wire flitsAreTail_5;
  wire T976;
  wire T977;
  wire T978;
  wire T979;
  wire[53:0] T980;
  wire T981;
  wire[30:0] T982;
  wire T983;
  wire T984;
  wire T985;
  wire T986;
  wire T987;
  wire[54:0] T988;
  wire[54:0] T989;
  wire T990;
  wire T991;
  wire T992;
  wire T993;
  wire T994;
  wire T995;
  wire T996;
  wire T997;
  wire T998;
  wire T999;
  wire[54:0] T1000;
  wire[54:0] T1001;
  wire T3147;
  reg [54:0] R1002;
  wire[54:0] T3148;
  wire[54:0] T1003;
  wire[54:0] T3149;
  wire T1004;
  wire T1005;
  wire[54:0] T1006;
  wire[54:0] T1007;
  wire T1008;
  wire T1009;
  wire[1:0] T1010;
  wire[1:0] T1011;
  wire[1:0] T1012;
  wire T1013;
  wire[2:0] T1014;
  reg [2:0] R1015;
  wire[2:0] T3150;
  wire[1:0] T1016;
  wire T1017;
  wire T1018;
  wire T1019;
  wire T1020;
  wire T1021;
  wire T1022;
  wire T1023;
  wire T1024;
  wire T1025;
  wire[2:0] T1026;
  wire T1027;
  wire T1028;
  wire T1029;
  wire T1030;
  wire T1031;
  wire T1032;
  wire T1033;
  wire T1034;
  wire T1035;
  wire T1036;
  wire T1037;
  wire T1038;
  wire T1039;
  wire T3151;
  wire T1040;
  wire T1041;
  wire[3:0] T1042;
  wire[3:0] T1043;
  wire[3:0] T1044;
  wire T1045;
  wire[2:0] T1046;
  wire[3:0] T1047;
  wire T1048;
  wire T1049;
  wire T1050;
  wire T1051;
  wire T1052;
  wire T1053;
  wire T1054;
  wire[2:0] T1055;
  wire T1056;
  wire T1057;
  wire T1058;
  wire T1059;
  wire T1060;
  wire T1061;
  wire T1062;
  wire T1063;
  wire[53:0] T1064;
  wire T1065;
  wire[30:0] T1066;
  wire T1067;
  wire T1068;
  reg  R1069;
  wire T3152;
  wire[2:0] T1070;
  wire[30:0] T1071;
  wire[54:0] T1072;
  wire[1:0] T1073;
  wire[1:0] T1074;
  wire[1:0] T1075;
  wire[3:0] T1076;
  wire T1077;
  wire T1078;
  wire[15:0] T1079;
  wire T1080;
  wire T1081;
  wire T1082;
  wire T1083;
  wire T1084;
  wire T1085;
  wire T1086;
  wire T1087;
  wire T1088;
  wire T1089;
  wire T1090;
  wire T1091;
  wire T1092;
  wire T1093;
  wire T1094;
  wire T1095;
  wire T1096;
  wire T1097;
  wire T1098;
  wire T1099;
  wire T1100;
  wire T1101;
  wire T1102;
  wire T1103;
  wire T1104;
  wire T1105;
  wire T1106;
  wire T1107;
  wire[54:0] T3153;
  wire[30:0] T1108;
  wire[30:0] T1109;
  wire[8:0] T1110;
  wire[4:0] T1111;
  wire[3:0] T1112;
  wire[21:0] T1113;
  wire[4:0] T1114;
  wire[16:0] T1115;
  wire T1116;
  wire T1117;
  wire T1118;
  wire T1119;
  wire flitsAreTail_4;
  wire T1120;
  wire T1121;
  wire T1122;
  wire T1123;
  wire[53:0] T1124;
  wire T1125;
  wire[30:0] T1126;
  wire T1127;
  wire T1128;
  wire T1129;
  wire T1130;
  wire T1131;
  wire[54:0] T1132;
  wire[54:0] T1133;
  wire T1134;
  wire T1135;
  wire T1136;
  wire T1137;
  wire T1138;
  wire T1139;
  wire T1140;
  wire T1141;
  wire T1142;
  wire T1143;
  wire[54:0] T1144;
  wire[54:0] T1145;
  wire T3154;
  reg [54:0] R1146;
  wire[54:0] T3155;
  wire[54:0] T1147;
  wire[54:0] T3156;
  wire T1148;
  wire T1149;
  wire[54:0] T1150;
  wire[54:0] T1151;
  wire T1152;
  wire T1153;
  wire[1:0] T1154;
  wire[1:0] T1155;
  wire[1:0] T1156;
  wire T1157;
  wire[2:0] T1158;
  reg [2:0] R1159;
  wire[2:0] T3157;
  wire[1:0] T1160;
  wire T1161;
  wire T1162;
  wire T1163;
  wire T1164;
  wire T1165;
  wire T1166;
  wire T1167;
  wire T1168;
  wire T1169;
  wire[2:0] T1170;
  wire T1171;
  wire T1172;
  wire T1173;
  wire T1174;
  wire T1175;
  wire T1176;
  wire T1177;
  wire T1178;
  wire T1179;
  wire T1180;
  wire T1181;
  wire T1182;
  wire T1183;
  wire T3158;
  wire T1184;
  wire T1185;
  wire[3:0] T1186;
  wire[3:0] T1187;
  wire[3:0] T1188;
  wire T1189;
  wire[2:0] T1190;
  wire[3:0] T1191;
  wire T1192;
  wire T1193;
  wire T1194;
  wire T1195;
  wire T1196;
  wire T1197;
  wire T1198;
  wire[2:0] T1199;
  wire T1200;
  wire T1201;
  wire T1202;
  wire T1203;
  wire T1204;
  wire T1205;
  wire T1206;
  wire T1207;
  wire[53:0] T1208;
  wire T1209;
  wire[30:0] T1210;
  wire T1211;
  wire T1212;
  reg  R1213;
  wire T3159;
  wire[2:0] T1214;
  wire[30:0] T1215;
  wire[54:0] T1216;
  wire[1:0] T1217;
  wire[1:0] T1218;
  wire[1:0] T1219;
  wire[3:0] T1220;
  wire T1221;
  wire T1222;
  wire[15:0] T1223;
  wire T1224;
  wire T1225;
  wire T1226;
  wire T1227;
  wire T1228;
  wire T1229;
  wire T1230;
  wire T1231;
  wire T1232;
  wire T1233;
  wire T1234;
  wire T1235;
  wire T1236;
  wire T1237;
  wire T1238;
  wire T1239;
  wire T1240;
  wire T1241;
  wire T1242;
  wire T1243;
  wire T1244;
  wire T1245;
  wire T1246;
  wire T1247;
  wire T1248;
  wire T1249;
  wire T1250;
  wire T1251;
  wire[54:0] T3160;
  wire[30:0] T1252;
  wire[30:0] T1253;
  wire[8:0] T1254;
  wire[4:0] T1255;
  wire[3:0] T1256;
  wire[21:0] T1257;
  wire[4:0] T1258;
  wire[16:0] T1259;
  wire T1260;
  wire T1261;
  wire T1262;
  wire T1263;
  wire flitsAreTail_3;
  wire T1264;
  wire T1265;
  wire T1266;
  wire T1267;
  wire[53:0] T1268;
  wire T1269;
  wire[30:0] T1270;
  wire T1271;
  wire T1272;
  wire T1273;
  wire T1274;
  wire T1275;
  wire[54:0] T1276;
  wire[54:0] T1277;
  wire T1278;
  wire T1279;
  wire T1280;
  wire T1281;
  wire T1282;
  wire T1283;
  wire T1284;
  wire T1285;
  wire T1286;
  wire T1287;
  wire[54:0] T1288;
  wire[54:0] T1289;
  wire T3161;
  reg [54:0] R1290;
  wire[54:0] T3162;
  wire[54:0] T1291;
  wire[54:0] T3163;
  wire T1292;
  wire T1293;
  wire[54:0] T1294;
  wire[54:0] T1295;
  wire T1296;
  wire T1297;
  wire[1:0] T1298;
  wire[1:0] T1299;
  wire[1:0] T1300;
  wire T1301;
  wire[2:0] T1302;
  reg [2:0] R1303;
  wire[2:0] T3164;
  wire[1:0] T1304;
  wire T1305;
  wire T1306;
  wire T1307;
  wire T1308;
  wire T1309;
  wire T1310;
  wire T1311;
  wire T1312;
  wire T1313;
  wire[2:0] T1314;
  wire T1315;
  wire T1316;
  wire T1317;
  wire T1318;
  wire T1319;
  wire T1320;
  wire T1321;
  wire T1322;
  wire T1323;
  wire T1324;
  wire T1325;
  wire T1326;
  wire T1327;
  wire T3165;
  wire T1328;
  wire T1329;
  wire[3:0] T1330;
  wire[3:0] T1331;
  wire[3:0] T1332;
  wire T1333;
  wire[2:0] T1334;
  wire[3:0] T1335;
  wire T1336;
  wire T1337;
  wire T1338;
  wire T1339;
  wire T1340;
  wire T1341;
  wire T1342;
  wire[2:0] T1343;
  wire T1344;
  wire T1345;
  wire T1346;
  wire T1347;
  wire T1348;
  wire T1349;
  wire T1350;
  wire T1351;
  wire[53:0] T1352;
  wire T1353;
  wire[30:0] T1354;
  wire T1355;
  wire T1356;
  reg  R1357;
  wire T3166;
  wire[2:0] T1358;
  wire[30:0] T1359;
  wire[54:0] T1360;
  wire[1:0] T1361;
  wire[1:0] T1362;
  wire[1:0] T1363;
  wire[3:0] T1364;
  wire T1365;
  wire T1366;
  wire[15:0] T1367;
  wire T1368;
  wire T1369;
  wire T1370;
  wire T1371;
  wire T1372;
  wire T1373;
  wire T1374;
  wire T1375;
  wire T1376;
  wire T1377;
  wire T1378;
  wire T1379;
  wire T1380;
  wire T1381;
  wire T1382;
  wire T1383;
  wire T1384;
  wire T1385;
  wire T1386;
  wire T1387;
  wire T1388;
  wire T1389;
  wire T1390;
  wire T1391;
  wire T1392;
  wire T1393;
  wire T1394;
  wire T1395;
  wire[54:0] T3167;
  wire[30:0] T1396;
  wire[30:0] T1397;
  wire[8:0] T1398;
  wire[4:0] T1399;
  wire[3:0] T1400;
  wire[21:0] T1401;
  wire[4:0] T1402;
  wire[16:0] T1403;
  wire T1404;
  wire T1405;
  wire T1406;
  wire T1407;
  wire flitsAreTail_2;
  wire T1408;
  wire T1409;
  wire T1410;
  wire T1411;
  wire[53:0] T1412;
  wire T1413;
  wire[30:0] T1414;
  wire T1415;
  wire T1416;
  wire T1417;
  wire T1418;
  wire T1419;
  wire[54:0] T1420;
  wire[54:0] T1421;
  wire T1422;
  wire T1423;
  wire T1424;
  wire T1425;
  wire T1426;
  wire T1427;
  wire T1428;
  wire T1429;
  wire T1430;
  wire T1431;
  wire[54:0] T1432;
  wire[54:0] T1433;
  wire T3168;
  reg [54:0] R1434;
  wire[54:0] T3169;
  wire[54:0] T1435;
  wire[54:0] T3170;
  wire T1436;
  wire T1437;
  wire[54:0] T1438;
  wire[54:0] T1439;
  wire T1440;
  wire T1441;
  wire[1:0] T1442;
  wire[1:0] T1443;
  wire[1:0] T1444;
  wire T1445;
  wire[2:0] T1446;
  reg [2:0] R1447;
  wire[2:0] T3171;
  wire[1:0] T1448;
  wire T1449;
  wire T1450;
  wire T1451;
  wire T1452;
  wire T1453;
  wire T1454;
  wire T1455;
  wire T1456;
  wire T1457;
  wire[2:0] T1458;
  wire T1459;
  wire T1460;
  wire T1461;
  wire T1462;
  wire T1463;
  wire T1464;
  wire T1465;
  wire T1466;
  wire T1467;
  wire T1468;
  wire T1469;
  wire T1470;
  wire T1471;
  wire T3172;
  wire T1472;
  wire T1473;
  wire[3:0] T1474;
  wire[3:0] T1475;
  wire[3:0] T1476;
  wire T1477;
  wire[2:0] T1478;
  wire[3:0] T1479;
  wire T1480;
  wire T1481;
  wire T1482;
  wire T1483;
  wire T1484;
  wire T1485;
  wire T1486;
  wire[2:0] T1487;
  wire T1488;
  wire T1489;
  wire T1490;
  wire T1491;
  wire T1492;
  wire T1493;
  wire T1494;
  wire T1495;
  wire[53:0] T1496;
  wire T1497;
  wire[30:0] T1498;
  wire T1499;
  wire T1500;
  reg  R1501;
  wire T3173;
  wire[2:0] T1502;
  wire[30:0] T1503;
  wire[54:0] T1504;
  wire[1:0] T1505;
  wire[1:0] T1506;
  wire[1:0] T1507;
  wire[3:0] T1508;
  wire T1509;
  wire T1510;
  wire[15:0] T1511;
  wire T1512;
  wire T1513;
  wire T1514;
  wire T1515;
  wire T1516;
  wire T1517;
  wire T1518;
  wire T1519;
  wire T1520;
  wire T1521;
  wire T1522;
  wire T1523;
  wire T1524;
  wire T1525;
  wire T1526;
  wire T1527;
  wire T1528;
  wire T1529;
  wire T1530;
  wire T1531;
  wire T1532;
  wire T1533;
  wire T1534;
  wire T1535;
  wire T1536;
  wire T1537;
  wire T1538;
  wire T1539;
  wire[54:0] T3174;
  wire[30:0] T1540;
  wire[30:0] T1541;
  wire[8:0] T1542;
  wire[4:0] T1543;
  wire[3:0] T1544;
  wire[21:0] T1545;
  wire[4:0] T1546;
  wire[16:0] T1547;
  wire T1548;
  wire T1549;
  wire T1550;
  wire T1551;
  wire flitsAreTail_1;
  wire T1552;
  wire T1553;
  wire T1554;
  wire T1555;
  wire[53:0] T1556;
  wire T1557;
  wire[30:0] T1558;
  wire T1559;
  wire T1560;
  wire T1561;
  wire T1562;
  wire T1563;
  wire[54:0] T1564;
  wire[54:0] T1565;
  wire T1566;
  wire T1567;
  wire T1568;
  wire T1569;
  wire T1570;
  wire T1571;
  wire T1572;
  wire T1573;
  wire T1574;
  wire T1575;
  wire[54:0] T1576;
  wire[54:0] T1577;
  wire T3175;
  reg [54:0] R1578;
  wire[54:0] T3176;
  wire[54:0] T1579;
  wire[54:0] T3177;
  wire T1580;
  wire T1581;
  wire[54:0] T1582;
  wire[54:0] T1583;
  wire T1584;
  wire T1585;
  wire[1:0] T1586;
  wire[1:0] T1587;
  wire[1:0] T1588;
  wire T1589;
  wire[2:0] T1590;
  reg [2:0] R1591;
  wire[2:0] T3178;
  wire[1:0] T1592;
  wire T1593;
  wire T1594;
  wire T1595;
  wire T1596;
  wire T1597;
  wire T1598;
  wire T1599;
  wire T1600;
  wire T1601;
  wire[2:0] T1602;
  wire T1603;
  wire T1604;
  wire T1605;
  wire T1606;
  wire T1607;
  wire T1608;
  wire T1609;
  wire T1610;
  wire T1611;
  wire T1612;
  wire T1613;
  wire T1614;
  wire T1615;
  wire T3179;
  wire T1616;
  wire T1617;
  wire[3:0] T1618;
  wire[3:0] T1619;
  wire[3:0] T1620;
  wire T1621;
  wire[2:0] T1622;
  wire[3:0] T1623;
  wire T1624;
  wire T1625;
  wire T1626;
  wire T1627;
  wire T1628;
  wire T1629;
  wire T1630;
  wire[2:0] T1631;
  wire T1632;
  wire T1633;
  wire T1634;
  wire T1635;
  wire T1636;
  wire T1637;
  wire T1638;
  wire T1639;
  wire[53:0] T1640;
  wire T1641;
  wire[30:0] T1642;
  wire T1643;
  wire T1644;
  reg  R1645;
  wire T3180;
  wire[2:0] T1646;
  wire[30:0] T1647;
  wire[54:0] T1648;
  wire[1:0] T1649;
  wire[1:0] T1650;
  wire[1:0] T1651;
  wire[3:0] T1652;
  wire T1653;
  wire T1654;
  wire[15:0] T1655;
  wire T1656;
  wire T1657;
  wire T1658;
  wire T1659;
  wire T1660;
  wire T1661;
  wire T1662;
  wire T1663;
  wire T1664;
  wire T1665;
  wire T1666;
  wire T1667;
  wire T1668;
  wire T1669;
  wire T1670;
  wire T1671;
  wire T1672;
  wire T1673;
  wire T1674;
  wire T1675;
  wire T1676;
  wire T1677;
  wire T1678;
  wire T1679;
  wire T1680;
  wire T1681;
  wire T1682;
  wire T1683;
  wire[54:0] T3181;
  wire[30:0] T1684;
  wire[30:0] T1685;
  wire[8:0] T1686;
  wire[4:0] T1687;
  wire[3:0] T1688;
  wire[21:0] T1689;
  wire[4:0] T1690;
  wire[16:0] T1691;
  wire T1692;
  wire T1693;
  wire T1694;
  wire T1695;
  wire flitsAreTail_0;
  wire T1696;
  wire T1697;
  wire T1698;
  wire T1699;
  wire[53:0] T1700;
  wire T1701;
  wire[30:0] T1702;
  wire T1703;
  wire T1704;
  wire T1705;
  wire T1706;
  wire T1707;
  wire[54:0] T1708;
  wire[54:0] T1709;
  wire T1710;
  wire T1711;
  wire T1712;
  wire T1713;
  wire T1714;
  wire T1715;
  wire T1716;
  wire T1717;
  wire T1718;
  wire T1719;
  wire T1720;
  wire T1721;
  wire T1722;
  wire[9:0] T1723;
  wire[9:0] T1724;
  wire[4:0] T1725;
  wire[2:0] T1726;
  wire[1:0] T1727;
  wire readyToXmit_0_4;
  wire T1728;
  wire T1729;
  wire T1730;
  wire T1731;
  wire T1732;
  wire T1733;
  wire T1734;
  wire T1735;
  wire[7:0] T1736;
  wire[2:0] T1737;
  wire T1738;
  wire T1739;
  wire T1740;
  wire T1741;
  wire T1742;
  wire T1743;
  wire T1744;
  wire readyToXmit_1_4;
  wire T1745;
  wire T1746;
  wire T1747;
  wire T1748;
  wire T1749;
  wire T1750;
  wire T1751;
  wire T1752;
  wire[7:0] T1753;
  wire[2:0] T1754;
  wire T1755;
  wire T1756;
  wire T1757;
  wire T1758;
  wire T1759;
  wire T1760;
  wire T1761;
  wire readyToXmit_2_4;
  wire T1762;
  wire T1763;
  wire T1764;
  wire T1765;
  wire T1766;
  wire T1767;
  wire T1768;
  wire T1769;
  wire[7:0] T1770;
  wire[2:0] T1771;
  wire T1772;
  wire T1773;
  wire T1774;
  wire T1775;
  wire T1776;
  wire T1777;
  wire T1778;
  wire[1:0] T1779;
  wire readyToXmit_3_4;
  wire T1780;
  wire T1781;
  wire T1782;
  wire T1783;
  wire T1784;
  wire T1785;
  wire T1786;
  wire T1787;
  wire[7:0] T1788;
  wire[2:0] T1789;
  wire T1790;
  wire T1791;
  wire T1792;
  wire T1793;
  wire T1794;
  wire T1795;
  wire T1796;
  wire readyToXmit_4_4;
  wire T1797;
  wire T1798;
  wire T1799;
  wire T1800;
  wire T1801;
  wire T1802;
  wire T1803;
  wire T1804;
  wire[7:0] T1805;
  wire[2:0] T1806;
  wire T1807;
  wire T1808;
  wire T1809;
  wire T1810;
  wire T1811;
  wire T1812;
  wire T1813;
  wire[4:0] T1814;
  wire[2:0] T1815;
  wire[1:0] T1816;
  wire readyToXmit_5_4;
  wire T1817;
  wire T1818;
  wire T1819;
  wire T1820;
  wire T1821;
  wire T1822;
  wire T1823;
  wire T1824;
  wire[7:0] T1825;
  wire[2:0] T1826;
  wire T1827;
  wire T1828;
  wire T1829;
  wire T1830;
  wire T1831;
  wire T1832;
  wire T1833;
  wire readyToXmit_6_4;
  wire T1834;
  wire T1835;
  wire T1836;
  wire T1837;
  wire T1838;
  wire T1839;
  wire T1840;
  wire T1841;
  wire[7:0] T1842;
  wire[2:0] T1843;
  wire T1844;
  wire T1845;
  wire T1846;
  wire T1847;
  wire T1848;
  wire T1849;
  wire T1850;
  wire readyToXmit_7_4;
  wire T1851;
  wire T1852;
  wire T1853;
  wire T1854;
  wire T1855;
  wire T1856;
  wire T1857;
  wire T1858;
  wire[7:0] T1859;
  wire[2:0] T1860;
  wire T1861;
  wire T1862;
  wire T1863;
  wire T1864;
  wire T1865;
  wire T1866;
  wire T1867;
  wire[1:0] T1868;
  wire readyToXmit_8_4;
  wire T1869;
  wire T1870;
  wire T1871;
  wire T1872;
  wire T1873;
  wire T1874;
  wire T1875;
  wire T1876;
  wire[7:0] T1877;
  wire[2:0] T1878;
  wire T1879;
  wire T1880;
  wire T1881;
  wire T1882;
  wire T1883;
  wire T1884;
  wire T1885;
  wire readyToXmit_9_4;
  wire T1886;
  wire T1887;
  wire T1888;
  wire T1889;
  wire T1890;
  wire T1891;
  wire T1892;
  wire T1893;
  wire[7:0] T1894;
  wire[2:0] T1895;
  wire T1896;
  wire T1897;
  wire T1898;
  wire T1899;
  wire T1900;
  wire T1901;
  wire T1902;
  wire T1903;
  wire T1904;
  wire T1905;
  wire[9:0] T1906;
  wire[9:0] T1907;
  wire[4:0] T1908;
  wire[2:0] T1909;
  wire[1:0] T1910;
  wire readyToXmit_0_3;
  wire T1911;
  wire T1912;
  wire T1913;
  wire T1914;
  wire T1915;
  wire readyToXmit_1_3;
  wire T1916;
  wire T1917;
  wire T1918;
  wire T1919;
  wire T1920;
  wire readyToXmit_2_3;
  wire T1921;
  wire T1922;
  wire T1923;
  wire T1924;
  wire T1925;
  wire[1:0] T1926;
  wire readyToXmit_3_3;
  wire T1927;
  wire T1928;
  wire T1929;
  wire T1930;
  wire T1931;
  wire readyToXmit_4_3;
  wire T1932;
  wire T1933;
  wire T1934;
  wire T1935;
  wire T1936;
  wire[4:0] T1937;
  wire[2:0] T1938;
  wire[1:0] T1939;
  wire readyToXmit_5_3;
  wire T1940;
  wire T1941;
  wire T1942;
  wire T1943;
  wire T1944;
  wire readyToXmit_6_3;
  wire T1945;
  wire T1946;
  wire T1947;
  wire T1948;
  wire T1949;
  wire readyToXmit_7_3;
  wire T1950;
  wire T1951;
  wire T1952;
  wire T1953;
  wire T1954;
  wire[1:0] T1955;
  wire readyToXmit_8_3;
  wire T1956;
  wire T1957;
  wire T1958;
  wire T1959;
  wire T1960;
  wire readyToXmit_9_3;
  wire T1961;
  wire T1962;
  wire T1963;
  wire T1964;
  wire T1965;
  wire T1966;
  wire T1967;
  wire T1968;
  wire[9:0] T1969;
  wire[9:0] T1970;
  wire[4:0] T1971;
  wire[2:0] T1972;
  wire[1:0] T1973;
  wire readyToXmit_0_2;
  wire T1974;
  wire T1975;
  wire T1976;
  wire T1977;
  wire T1978;
  wire readyToXmit_1_2;
  wire T1979;
  wire T1980;
  wire T1981;
  wire T1982;
  wire T1983;
  wire readyToXmit_2_2;
  wire T1984;
  wire T1985;
  wire T1986;
  wire T1987;
  wire T1988;
  wire[1:0] T1989;
  wire readyToXmit_3_2;
  wire T1990;
  wire T1991;
  wire T1992;
  wire T1993;
  wire T1994;
  wire readyToXmit_4_2;
  wire T1995;
  wire T1996;
  wire T1997;
  wire T1998;
  wire T1999;
  wire[4:0] T2000;
  wire[2:0] T2001;
  wire[1:0] T2002;
  wire readyToXmit_5_2;
  wire T2003;
  wire T2004;
  wire T2005;
  wire T2006;
  wire T2007;
  wire readyToXmit_6_2;
  wire T2008;
  wire T2009;
  wire T2010;
  wire T2011;
  wire T2012;
  wire readyToXmit_7_2;
  wire T2013;
  wire T2014;
  wire T2015;
  wire T2016;
  wire T2017;
  wire[1:0] T2018;
  wire readyToXmit_8_2;
  wire T2019;
  wire T2020;
  wire T2021;
  wire T2022;
  wire T2023;
  wire readyToXmit_9_2;
  wire T2024;
  wire T2025;
  wire T2026;
  wire T2027;
  wire T2028;
  wire T2029;
  wire T2030;
  wire T2031;
  wire[9:0] T2032;
  wire[9:0] T2033;
  wire[4:0] T2034;
  wire[2:0] T2035;
  wire[1:0] T2036;
  wire readyToXmit_0_1;
  wire T2037;
  wire T2038;
  wire T2039;
  wire T2040;
  wire T2041;
  wire readyToXmit_1_1;
  wire T2042;
  wire T2043;
  wire T2044;
  wire T2045;
  wire T2046;
  wire readyToXmit_2_1;
  wire T2047;
  wire T2048;
  wire T2049;
  wire T2050;
  wire T2051;
  wire[1:0] T2052;
  wire readyToXmit_3_1;
  wire T2053;
  wire T2054;
  wire T2055;
  wire T2056;
  wire T2057;
  wire readyToXmit_4_1;
  wire T2058;
  wire T2059;
  wire T2060;
  wire T2061;
  wire T2062;
  wire[4:0] T2063;
  wire[2:0] T2064;
  wire[1:0] T2065;
  wire readyToXmit_5_1;
  wire T2066;
  wire T2067;
  wire T2068;
  wire T2069;
  wire T2070;
  wire readyToXmit_6_1;
  wire T2071;
  wire T2072;
  wire T2073;
  wire T2074;
  wire T2075;
  wire readyToXmit_7_1;
  wire T2076;
  wire T2077;
  wire T2078;
  wire T2079;
  wire T2080;
  wire[1:0] T2081;
  wire readyToXmit_8_1;
  wire T2082;
  wire T2083;
  wire T2084;
  wire T2085;
  wire T2086;
  wire readyToXmit_9_1;
  wire T2087;
  wire T2088;
  wire T2089;
  wire T2090;
  wire T2091;
  wire T2092;
  wire T2093;
  wire T2094;
  wire[9:0] T2095;
  wire[9:0] T2096;
  wire[4:0] T2097;
  wire[2:0] T2098;
  wire[1:0] T2099;
  wire readyToXmit_0_0;
  wire T2100;
  wire T2101;
  wire T2102;
  wire T2103;
  wire T2104;
  wire readyToXmit_1_0;
  wire T2105;
  wire T2106;
  wire T2107;
  wire T2108;
  wire T2109;
  wire readyToXmit_2_0;
  wire T2110;
  wire T2111;
  wire T2112;
  wire T2113;
  wire T2114;
  wire[1:0] T2115;
  wire readyToXmit_3_0;
  wire T2116;
  wire T2117;
  wire T2118;
  wire T2119;
  wire T2120;
  wire readyToXmit_4_0;
  wire T2121;
  wire T2122;
  wire T2123;
  wire T2124;
  wire T2125;
  wire[4:0] T2126;
  wire[2:0] T2127;
  wire[1:0] T2128;
  wire readyToXmit_5_0;
  wire T2129;
  wire T2130;
  wire T2131;
  wire T2132;
  wire T2133;
  wire readyToXmit_6_0;
  wire T2134;
  wire T2135;
  wire T2136;
  wire T2137;
  wire T2138;
  wire readyToXmit_7_0;
  wire T2139;
  wire T2140;
  wire T2141;
  wire T2142;
  wire T2143;
  wire[1:0] T2144;
  wire readyToXmit_8_0;
  wire T2145;
  wire T2146;
  wire T2147;
  wire T2148;
  wire T2149;
  wire readyToXmit_9_0;
  wire T2150;
  wire T2151;
  wire T2152;
  wire T2153;
  wire T2154;
  wire T2155;
  wire T2156;
  wire T2157;
  wire T2158;
  wire T2159;
  wire T2160;
  wire T2161;
  wire T2162;
  wire T2163;
  wire T2164;
  wire T2165;
  wire T2166;
  wire T2167;
  wire T2168;
  wire T2169;
  wire T2170;
  wire T2171;
  wire T2172;
  wire T2173;
  wire T2174;
  wire T2175;
  reg [1:0] validVCs_0_0;
  reg  R2176;
  wire T2177;
  wire T2178;
  wire T2179;
  wire T2180;
  reg  R2181;
  wire T2182;
  wire T2183;
  wire T2184;
  wire T2185;
  reg [1:0] validVCs_0_1;
  reg  R2186;
  wire T2187;
  wire T2188;
  wire T2189;
  wire T2190;
  reg  R2191;
  wire T2192;
  wire T2193;
  wire T2194;
  wire T2195;
  reg [1:0] validVCs_0_2;
  reg  R2196;
  wire T2197;
  wire T2198;
  wire T2199;
  wire T2200;
  reg  R2201;
  wire T2202;
  wire T2203;
  wire T2204;
  wire T2205;
  reg [1:0] validVCs_0_3;
  reg  R2206;
  wire T2207;
  wire T2208;
  wire T2209;
  wire T2210;
  reg  R2211;
  wire T2212;
  wire T2213;
  wire T2214;
  wire T2215;
  reg [1:0] validVCs_0_4;
  reg  R2216;
  wire T2217;
  wire T2218;
  wire T2219;
  wire T2220;
  reg  R2221;
  wire T2222;
  wire T2223;
  wire T2224;
  wire T2225;
  reg [1:0] validVCs_1_0;
  reg  R2226;
  wire T2227;
  wire T2228;
  wire T2229;
  wire T2230;
  reg  R2231;
  wire T2232;
  wire T2233;
  wire T2234;
  wire T2235;
  reg [1:0] validVCs_1_1;
  reg  R2236;
  wire T2237;
  wire T2238;
  wire T2239;
  wire T2240;
  reg  R2241;
  wire T2242;
  wire T2243;
  wire T2244;
  wire T2245;
  reg [1:0] validVCs_1_2;
  reg  R2246;
  wire T2247;
  wire T2248;
  wire T2249;
  wire T2250;
  reg  R2251;
  wire T2252;
  wire T2253;
  wire T2254;
  wire T2255;
  reg [1:0] validVCs_1_3;
  reg  R2256;
  wire T2257;
  wire T2258;
  wire T2259;
  wire T2260;
  reg  R2261;
  wire T2262;
  wire T2263;
  wire T2264;
  wire T2265;
  reg [1:0] validVCs_1_4;
  reg  R2266;
  wire T2267;
  wire T2268;
  wire T2269;
  wire T2270;
  reg  R2271;
  wire T2272;
  wire T2273;
  wire T2274;
  wire T2275;
  reg [1:0] validVCs_2_0;
  reg  R2276;
  wire T2277;
  wire T2278;
  wire T2279;
  wire T2280;
  reg  R2281;
  wire T2282;
  wire T2283;
  wire T2284;
  wire T2285;
  reg [1:0] validVCs_2_1;
  reg  R2286;
  wire T2287;
  wire T2288;
  wire T2289;
  wire T2290;
  reg  R2291;
  wire T2292;
  wire T2293;
  wire T2294;
  wire T2295;
  reg [1:0] validVCs_2_2;
  reg  R2296;
  wire T2297;
  wire T2298;
  wire T2299;
  wire T2300;
  reg  R2301;
  wire T2302;
  wire T2303;
  wire T2304;
  wire T2305;
  reg [1:0] validVCs_2_3;
  reg  R2306;
  wire T2307;
  wire T2308;
  wire T2309;
  wire T2310;
  reg  R2311;
  wire T2312;
  wire T2313;
  wire T2314;
  wire T2315;
  reg [1:0] validVCs_2_4;
  reg  R2316;
  wire T2317;
  wire T2318;
  wire T2319;
  wire T2320;
  reg  R2321;
  wire T2322;
  wire T2323;
  wire T2324;
  wire T2325;
  reg [1:0] validVCs_3_0;
  reg  R2326;
  wire T2327;
  wire T2328;
  wire T2329;
  wire T2330;
  reg  R2331;
  wire T2332;
  wire T2333;
  wire T2334;
  wire T2335;
  reg [1:0] validVCs_3_1;
  reg  R2336;
  wire T2337;
  wire T2338;
  wire T2339;
  wire T2340;
  reg  R2341;
  wire T2342;
  wire T2343;
  wire T2344;
  wire T2345;
  reg [1:0] validVCs_3_2;
  reg  R2346;
  wire T2347;
  wire T2348;
  wire T2349;
  wire T2350;
  reg  R2351;
  wire T2352;
  wire T2353;
  wire T2354;
  wire T2355;
  reg [1:0] validVCs_3_3;
  reg  R2356;
  wire T2357;
  wire T2358;
  wire T2359;
  wire T2360;
  reg  R2361;
  wire T2362;
  wire T2363;
  wire T2364;
  wire T2365;
  reg [1:0] validVCs_3_4;
  reg  R2366;
  wire T2367;
  wire T2368;
  wire T2369;
  wire T2370;
  reg  R2371;
  wire T2372;
  wire T2373;
  wire T2374;
  wire T2375;
  reg [1:0] validVCs_4_0;
  reg  R2376;
  wire T2377;
  wire T2378;
  wire T2379;
  wire T2380;
  reg  R2381;
  wire T2382;
  wire T2383;
  wire T2384;
  wire T2385;
  reg [1:0] validVCs_4_1;
  reg  R2386;
  wire T2387;
  wire T2388;
  wire T2389;
  wire T2390;
  reg  R2391;
  wire T2392;
  wire T2393;
  wire T2394;
  wire T2395;
  reg [1:0] validVCs_4_2;
  reg  R2396;
  wire T2397;
  wire T2398;
  wire T2399;
  wire T2400;
  reg  R2401;
  wire T2402;
  wire T2403;
  wire T2404;
  wire T2405;
  reg [1:0] validVCs_4_3;
  reg  R2406;
  wire T2407;
  wire T2408;
  wire T2409;
  wire T2410;
  reg  R2411;
  wire T2412;
  wire T2413;
  wire T2414;
  wire T2415;
  reg [1:0] validVCs_4_4;
  reg  R2416;
  wire T2417;
  wire T2418;
  wire T2419;
  wire T2420;
  reg  R2421;
  wire T2422;
  wire T2423;
  wire T2424;
  wire T2425;
  reg [1:0] validVCs_5_0;
  reg  R2426;
  wire T2427;
  wire T2428;
  wire T2429;
  wire T2430;
  reg  R2431;
  wire T2432;
  wire T2433;
  wire T2434;
  wire T2435;
  reg [1:0] validVCs_5_1;
  reg  R2436;
  wire T2437;
  wire T2438;
  wire T2439;
  wire T2440;
  reg  R2441;
  wire T2442;
  wire T2443;
  wire T2444;
  wire T2445;
  reg [1:0] validVCs_5_2;
  reg  R2446;
  wire T2447;
  wire T2448;
  wire T2449;
  wire T2450;
  reg  R2451;
  wire T2452;
  wire T2453;
  wire T2454;
  wire T2455;
  reg [1:0] validVCs_5_3;
  reg  R2456;
  wire T2457;
  wire T2458;
  wire T2459;
  wire T2460;
  reg  R2461;
  wire T2462;
  wire T2463;
  wire T2464;
  wire T2465;
  reg [1:0] validVCs_5_4;
  reg  R2466;
  wire T2467;
  wire T2468;
  wire T2469;
  wire T2470;
  reg  R2471;
  wire T2472;
  wire T2473;
  wire T2474;
  wire T2475;
  reg [1:0] validVCs_6_0;
  reg  R2476;
  wire T2477;
  wire T2478;
  wire T2479;
  wire T2480;
  reg  R2481;
  wire T2482;
  wire T2483;
  wire T2484;
  wire T2485;
  reg [1:0] validVCs_6_1;
  reg  R2486;
  wire T2487;
  wire T2488;
  wire T2489;
  wire T2490;
  reg  R2491;
  wire T2492;
  wire T2493;
  wire T2494;
  wire T2495;
  reg [1:0] validVCs_6_2;
  reg  R2496;
  wire T2497;
  wire T2498;
  wire T2499;
  wire T2500;
  reg  R2501;
  wire T2502;
  wire T2503;
  wire T2504;
  wire T2505;
  reg [1:0] validVCs_6_3;
  reg  R2506;
  wire T2507;
  wire T2508;
  wire T2509;
  wire T2510;
  reg  R2511;
  wire T2512;
  wire T2513;
  wire T2514;
  wire T2515;
  reg [1:0] validVCs_6_4;
  reg  R2516;
  wire T2517;
  wire T2518;
  wire T2519;
  wire T2520;
  reg  R2521;
  wire T2522;
  wire T2523;
  wire T2524;
  wire T2525;
  reg [1:0] validVCs_7_0;
  reg  R2526;
  wire T2527;
  wire T2528;
  wire T2529;
  wire T2530;
  reg  R2531;
  wire T2532;
  wire T2533;
  wire T2534;
  wire T2535;
  reg [1:0] validVCs_7_1;
  reg  R2536;
  wire T2537;
  wire T2538;
  wire T2539;
  wire T2540;
  reg  R2541;
  wire T2542;
  wire T2543;
  wire T2544;
  wire T2545;
  reg [1:0] validVCs_7_2;
  reg  R2546;
  wire T2547;
  wire T2548;
  wire T2549;
  wire T2550;
  reg  R2551;
  wire T2552;
  wire T2553;
  wire T2554;
  wire T2555;
  reg [1:0] validVCs_7_3;
  reg  R2556;
  wire T2557;
  wire T2558;
  wire T2559;
  wire T2560;
  reg  R2561;
  wire T2562;
  wire T2563;
  wire T2564;
  wire T2565;
  reg [1:0] validVCs_7_4;
  reg  R2566;
  wire T2567;
  wire T2568;
  wire T2569;
  wire T2570;
  reg  R2571;
  wire T2572;
  wire T2573;
  wire T2574;
  wire T2575;
  reg [1:0] validVCs_8_0;
  reg  R2576;
  wire T2577;
  wire T2578;
  wire T2579;
  wire T2580;
  reg  R2581;
  wire T2582;
  wire T2583;
  wire T2584;
  wire T2585;
  reg [1:0] validVCs_8_1;
  reg  R2586;
  wire T2587;
  wire T2588;
  wire T2589;
  wire T2590;
  reg  R2591;
  wire T2592;
  wire T2593;
  wire T2594;
  wire T2595;
  reg [1:0] validVCs_8_2;
  reg  R2596;
  wire T2597;
  wire T2598;
  wire T2599;
  wire T2600;
  reg  R2601;
  wire T2602;
  wire T2603;
  wire T2604;
  wire T2605;
  reg [1:0] validVCs_8_3;
  reg  R2606;
  wire T2607;
  wire T2608;
  wire T2609;
  wire T2610;
  reg  R2611;
  wire T2612;
  wire T2613;
  wire T2614;
  wire T2615;
  reg [1:0] validVCs_8_4;
  reg  R2616;
  wire T2617;
  wire T2618;
  wire T2619;
  wire T2620;
  reg  R2621;
  wire T2622;
  wire T2623;
  wire T2624;
  wire T2625;
  reg [1:0] validVCs_9_0;
  reg  R2626;
  wire T2627;
  wire T2628;
  wire T2629;
  wire T2630;
  reg  R2631;
  wire T2632;
  wire T2633;
  wire T2634;
  wire T2635;
  reg [1:0] validVCs_9_1;
  reg  R2636;
  wire T2637;
  wire T2638;
  wire T2639;
  wire T2640;
  reg  R2641;
  wire T2642;
  wire T2643;
  wire T2644;
  wire T2645;
  reg [1:0] validVCs_9_2;
  reg  R2646;
  wire T2647;
  wire T2648;
  wire T2649;
  wire T2650;
  reg  R2651;
  wire T2652;
  wire T2653;
  wire T2654;
  wire T2655;
  reg [1:0] validVCs_9_3;
  reg  R2656;
  wire T2657;
  wire T2658;
  wire T2659;
  wire T2660;
  reg  R2661;
  wire T2662;
  wire T2663;
  wire T2664;
  wire T2665;
  reg [1:0] validVCs_9_4;
  reg  R2666;
  wire T2667;
  wire T2668;
  wire T2669;
  wire T2670;
  reg  R2671;
  wire T2672;
  wire T2673;
  wire T2674;
  reg [2:0] R2675;
  wire[2:0] T3182;
  wire[2:0] T2676;
  wire[2:0] T2677;
  wire[30:0] T2678;
  wire T2679;
  wire T2680;
  wire T2681;
  wire T2682;
  reg [7:0] R2683;
  wire[7:0] T3183;
  wire[7:0] T2684;
  wire T2685;
  wire T2686;
  wire T2687;
  reg  R2688;
  wire T3184;
  reg [2:0] R2689;
  wire[2:0] T3185;
  wire[2:0] T2690;
  wire[2:0] T2691;
  wire[30:0] T2692;
  wire T2693;
  wire T2694;
  wire T2695;
  wire T2696;
  reg [7:0] R2697;
  wire[7:0] T3186;
  wire[7:0] T2698;
  wire T2699;
  wire T2700;
  wire T2701;
  reg  R2702;
  wire T3187;
  reg [2:0] R2703;
  wire[2:0] T3188;
  wire[2:0] T2704;
  wire[2:0] T2705;
  wire[30:0] T2706;
  wire T2707;
  wire T2708;
  wire T2709;
  wire T2710;
  reg [7:0] R2711;
  wire[7:0] T3189;
  wire[7:0] T2712;
  wire T2713;
  wire T2714;
  wire T2715;
  reg  R2716;
  wire T3190;
  reg [2:0] R2717;
  wire[2:0] T3191;
  wire[2:0] T2718;
  wire[2:0] T2719;
  wire[30:0] T2720;
  wire T2721;
  wire T2722;
  wire T2723;
  wire T2724;
  reg [7:0] R2725;
  wire[7:0] T3192;
  wire[7:0] T2726;
  wire T2727;
  wire T2728;
  wire T2729;
  reg  R2730;
  wire T3193;
  reg [2:0] R2731;
  wire[2:0] T3194;
  wire[2:0] T2732;
  wire[2:0] T2733;
  wire[30:0] T2734;
  wire T2735;
  wire T2736;
  wire T2737;
  wire T2738;
  reg [7:0] R2739;
  wire[7:0] T3195;
  wire[7:0] T2740;
  wire T2741;
  wire T2742;
  wire T2743;
  reg  R2744;
  wire T3196;
  reg [2:0] R2745;
  wire[2:0] T3197;
  wire[2:0] T2746;
  wire[2:0] T2747;
  wire[30:0] T2748;
  wire T2749;
  wire T2750;
  wire T2751;
  wire T2752;
  reg [7:0] R2753;
  wire[7:0] T3198;
  wire[7:0] T2754;
  wire T2755;
  wire T2756;
  wire T2757;
  reg  R2758;
  wire T3199;
  reg [2:0] R2759;
  wire[2:0] T3200;
  wire[2:0] T2760;
  wire[2:0] T2761;
  wire[30:0] T2762;
  wire T2763;
  wire T2764;
  wire T2765;
  wire T2766;
  reg [7:0] R2767;
  wire[7:0] T3201;
  wire[7:0] T2768;
  wire T2769;
  wire T2770;
  wire T2771;
  reg  R2772;
  wire T3202;
  reg [2:0] R2773;
  wire[2:0] T3203;
  wire[2:0] T2774;
  wire[2:0] T2775;
  wire[30:0] T2776;
  wire T2777;
  wire T2778;
  wire T2779;
  wire T2780;
  reg [7:0] R2781;
  wire[7:0] T3204;
  wire[7:0] T2782;
  wire T2783;
  wire T2784;
  wire T2785;
  reg  R2786;
  wire T3205;
  reg [2:0] R2787;
  wire[2:0] T3206;
  wire[2:0] T2788;
  wire[2:0] T2789;
  wire[30:0] T2790;
  wire T2791;
  wire T2792;
  wire T2793;
  wire T2794;
  reg [7:0] R2795;
  wire[7:0] T3207;
  wire[7:0] T2796;
  wire T2797;
  wire T2798;
  wire T2799;
  reg  R2800;
  wire T3208;
  reg [2:0] R2801;
  wire[2:0] T3209;
  wire[2:0] T2802;
  wire[2:0] T2803;
  wire[30:0] T2804;
  wire T2805;
  wire T2806;
  wire T2807;
  wire T2808;
  reg [7:0] R2809;
  wire[7:0] T3210;
  wire[7:0] T2810;
  wire T2811;
  wire T2812;
  wire T2813;
  reg  R2814;
  wire T3211;
  wire T2815;
  wire T2816;
  wire T2817;
  wire T2818;
  wire T2819;
  wire T2820;
  wire T2821;
  wire T2822;
  wire T2823;
  wire T2824;
  wire T2825;
  wire T2826;
  wire T2827;
  wire T2828;
  wire T2829;
  wire T2830;
  wire T2831;
  wire T2832;
  wire T2833;
  wire T2834;
  wire T2835;
  wire T2836;
  wire T2837;
  wire T2838;
  wire T2839;
  wire T2840;
  wire T2841;
  wire T2842;
  wire T2843;
  wire T2844;
  wire T2845;
  wire T2846;
  wire T2847;
  wire T2848;
  wire T2849;
  wire T2850;
  wire T2851;
  wire T2852;
  wire T2853;
  wire T2854;
  wire T2855;
  wire T2856;
  wire T2857;
  wire T2858;
  wire T2859;
  wire T2860;
  wire T2861;
  wire T2862;
  wire T2863;
  wire T2864;
  wire T2865;
  wire T2866;
  wire T2867;
  wire T2868;
  wire T2869;
  wire T2870;
  wire T2871;
  wire T2872;
  wire T2873;
  wire T2874;
  wire T2875;
  wire T2876;
  wire T2877;
  wire T2878;
  wire T2879;
  wire T2880;
  wire T2881;
  wire T2882;
  wire T2883;
  wire T2884;
  wire T2885;
  wire T2886;
  wire T2887;
  wire T2888;
  wire T2889;
  wire T2890;
  wire T2891;
  wire T2892;
  wire T2893;
  wire T2894;
  wire T2895;
  wire T2896;
  wire T2897;
  wire T2898;
  wire T2899;
  wire T2900;
  wire T2901;
  wire T2902;
  wire T2903;
  wire T2904;
  wire T2905;
  wire T2906;
  wire T2907;
  wire T2908;
  wire T2909;
  wire T2910;
  wire T2911;
  wire T2912;
  wire T2913;
  wire T2914;
  wire T2915;
  wire T2916;
  wire T2917;
  wire T2918;
  wire T2919;
  wire T2920;
  wire T2921;
  wire T2922;
  wire T2923;
  wire T2924;
  wire T2925;
  wire T2926;
  wire T2927;
  wire T2928;
  wire T2929;
  wire T2930;
  wire T2931;
  wire T2932;
  wire T2933;
  wire T2934;
  wire T2935;
  wire T2936;
  wire T2937;
  wire T2938;
  wire T2939;
  wire T2940;
  wire T2941;
  wire T2942;
  wire T2943;
  wire T2944;
  wire T2945;
  wire T2946;
  wire T2947;
  wire T2948;
  wire T2949;
  wire T2950;
  wire T2951;
  wire T2952;
  wire T2953;
  wire T2954;
  wire T2955;
  wire T2956;
  wire T2957;
  wire T2958;
  wire T2959;
  wire T2960;
  wire T2961;
  wire T2962;
  wire T2963;
  wire T2964;
  wire T2965;
  wire T2966;
  wire T2967;
  wire T2968;
  wire T2969;
  wire T2970;
  wire T2971;
  wire T2972;
  wire T2973;
  wire T2974;
  wire T2975;
  wire T2976;
  wire T2977;
  wire T2978;
  wire T2979;
  wire T2980;
  wire T2981;
  wire T2982;
  wire T2983;
  wire T2984;
  wire T2985;
  wire T2986;
  wire T2987;
  wire T2988;
  wire T2989;
  wire T2990;
  wire T2991;
  wire T2992;
  wire T2993;
  wire T2994;
  wire T2995;
  wire T2996;
  wire T2997;
  wire T2998;
  wire T2999;
  wire T3000;
  wire T3001;
  wire T3002;
  wire T3003;
  wire T3004;
  wire T3005;
  wire T3006;
  wire T3007;
  wire T3008;
  wire T3009;
  wire T3010;
  wire T3011;
  wire T3012;
  wire T3013;
  wire T3014;
  wire T3015;
  wire T3016;
  wire T3017;
  wire T3018;
  wire T3019;
  wire T3020;
  wire T3021;
  wire T3022;
  wire T3023;
  wire T3024;
  wire T3025;
  wire T3026;
  wire T3027;
  wire T3028;
  wire T3029;
  wire T3030;
  wire T3031;
  wire T3032;
  wire T3033;
  wire T3034;
  wire T3035;
  wire T3036;
  wire T3037;
  wire T3038;
  wire T3039;
  wire T3040;
  wire T3041;
  wire T3042;
  wire T3043;
  wire T3044;
  wire T3045;
  wire T3046;
  wire T3047;
  wire T3048;
  wire T3049;
  wire T3050;
  wire T3051;
  wire T3052;
  wire T3053;
  wire T3054;
  wire T3055;
  wire T3056;
  wire T3057;
  wire T3058;
  wire T3059;
  wire T3060;
  wire T3061;
  wire T3062;
  wire T3063;
  wire T3064;
  wire T3065;
  wire T3066;
  wire T3067;
  wire T3068;
  wire T3069;
  wire T3070;
  wire T3071;
  wire T3072;
  wire T3073;
  wire T3074;
  wire T3075;
  wire T3076;
  wire T3077;
  wire T3078;
  wire T3079;
  wire T3080;
  wire T3081;
  wire T3082;
  wire T3083;
  wire T3084;
  wire T3085;
  wire T3086;
  wire T3087;
  wire T3088;
  wire T3089;
  wire T3090;
  wire T3091;
  wire T3092;
  wire T3093;
  wire T3094;
  wire[31:0] T3212;
  wire T3095;
  wire T3096;
  reg  R3097;
  reg [54:0] R3098;
  wire[54:0] T3099;
  wire[54:0] T3213;
  reg  R3100;
  reg [54:0] R3101;
  wire[54:0] T3102;
  wire[54:0] T3214;
  reg  R3103;
  reg [54:0] R3104;
  wire[54:0] T3105;
  wire[54:0] T3215;
  reg  R3106;
  reg [54:0] R3107;
  wire[54:0] T3108;
  wire[54:0] T3216;
  reg  R3109;
  reg [54:0] R3110;
  wire[54:0] T3111;
  wire[54:0] T3217;
  wire[1:0] VCRouterOutputStateManagement_io_currentState;
  wire[1:0] VCRouterOutputStateManagement_1_io_currentState;
  wire[1:0] VCRouterOutputStateManagement_2_io_currentState;
  wire[1:0] VCRouterOutputStateManagement_3_io_currentState;
  wire[1:0] VCRouterOutputStateManagement_4_io_currentState;
  wire CreditGen_io_outCredit_grant;
  wire[54:0] RouterRegFile_io_readData;
  wire RouterRegFile_io_readValid;
  wire[54:0] RouterRegFile_io_readPipelineReg_1;
  wire[54:0] RouterRegFile_io_readPipelineReg_0;
  wire RouterRegFile_io_rvPipelineReg_1;
  wire RouterRegFile_io_rvPipelineReg_0;
  wire[15:0] CMeshDOR_io_outHeadFlit_packetID;
  wire CMeshDOR_io_outHeadFlit_isTail;
  wire CMeshDOR_io_outHeadFlit_vcPort;
  wire[3:0] CMeshDOR_io_outHeadFlit_packetType;
  wire[1:0] CMeshDOR_io_outHeadFlit_destination_2;
  wire[1:0] CMeshDOR_io_outHeadFlit_destination_1;
  wire[1:0] CMeshDOR_io_outHeadFlit_destination_0;
  wire[2:0] CMeshDOR_io_outHeadFlit_priorityLevel;
  wire[2:0] CMeshDOR_io_result;
  wire[1:0] CMeshDOR_io_vcsAvailable_4;
  wire[1:0] CMeshDOR_io_vcsAvailable_3;
  wire[1:0] CMeshDOR_io_vcsAvailable_2;
  wire[1:0] CMeshDOR_io_vcsAvailable_1;
  wire[1:0] CMeshDOR_io_vcsAvailable_0;
  wire[2:0] VCRouterStateManagement_io_currentState;
  wire CreditGen_1_io_outCredit_grant;
  wire[54:0] RouterRegFile_1_io_readData;
  wire RouterRegFile_1_io_readValid;
  wire[54:0] RouterRegFile_1_io_readPipelineReg_1;
  wire[54:0] RouterRegFile_1_io_readPipelineReg_0;
  wire RouterRegFile_1_io_rvPipelineReg_1;
  wire RouterRegFile_1_io_rvPipelineReg_0;
  wire[15:0] CMeshDOR_1_io_outHeadFlit_packetID;
  wire CMeshDOR_1_io_outHeadFlit_isTail;
  wire CMeshDOR_1_io_outHeadFlit_vcPort;
  wire[3:0] CMeshDOR_1_io_outHeadFlit_packetType;
  wire[1:0] CMeshDOR_1_io_outHeadFlit_destination_2;
  wire[1:0] CMeshDOR_1_io_outHeadFlit_destination_1;
  wire[1:0] CMeshDOR_1_io_outHeadFlit_destination_0;
  wire[2:0] CMeshDOR_1_io_outHeadFlit_priorityLevel;
  wire[2:0] CMeshDOR_1_io_result;
  wire[1:0] CMeshDOR_1_io_vcsAvailable_4;
  wire[1:0] CMeshDOR_1_io_vcsAvailable_3;
  wire[1:0] CMeshDOR_1_io_vcsAvailable_2;
  wire[1:0] CMeshDOR_1_io_vcsAvailable_1;
  wire[1:0] CMeshDOR_1_io_vcsAvailable_0;
  wire[2:0] VCRouterStateManagement_1_io_currentState;
  wire CreditGen_2_io_outCredit_grant;
  wire[54:0] RouterRegFile_2_io_readData;
  wire RouterRegFile_2_io_readValid;
  wire[54:0] RouterRegFile_2_io_readPipelineReg_1;
  wire[54:0] RouterRegFile_2_io_readPipelineReg_0;
  wire RouterRegFile_2_io_rvPipelineReg_1;
  wire RouterRegFile_2_io_rvPipelineReg_0;
  wire[15:0] CMeshDOR_2_io_outHeadFlit_packetID;
  wire CMeshDOR_2_io_outHeadFlit_isTail;
  wire CMeshDOR_2_io_outHeadFlit_vcPort;
  wire[3:0] CMeshDOR_2_io_outHeadFlit_packetType;
  wire[1:0] CMeshDOR_2_io_outHeadFlit_destination_2;
  wire[1:0] CMeshDOR_2_io_outHeadFlit_destination_1;
  wire[1:0] CMeshDOR_2_io_outHeadFlit_destination_0;
  wire[2:0] CMeshDOR_2_io_outHeadFlit_priorityLevel;
  wire[2:0] CMeshDOR_2_io_result;
  wire[1:0] CMeshDOR_2_io_vcsAvailable_4;
  wire[1:0] CMeshDOR_2_io_vcsAvailable_3;
  wire[1:0] CMeshDOR_2_io_vcsAvailable_2;
  wire[1:0] CMeshDOR_2_io_vcsAvailable_1;
  wire[1:0] CMeshDOR_2_io_vcsAvailable_0;
  wire[2:0] VCRouterStateManagement_2_io_currentState;
  wire CreditGen_3_io_outCredit_grant;
  wire[54:0] RouterRegFile_3_io_readData;
  wire RouterRegFile_3_io_readValid;
  wire[54:0] RouterRegFile_3_io_readPipelineReg_1;
  wire[54:0] RouterRegFile_3_io_readPipelineReg_0;
  wire RouterRegFile_3_io_rvPipelineReg_1;
  wire RouterRegFile_3_io_rvPipelineReg_0;
  wire[15:0] CMeshDOR_3_io_outHeadFlit_packetID;
  wire CMeshDOR_3_io_outHeadFlit_isTail;
  wire CMeshDOR_3_io_outHeadFlit_vcPort;
  wire[3:0] CMeshDOR_3_io_outHeadFlit_packetType;
  wire[1:0] CMeshDOR_3_io_outHeadFlit_destination_2;
  wire[1:0] CMeshDOR_3_io_outHeadFlit_destination_1;
  wire[1:0] CMeshDOR_3_io_outHeadFlit_destination_0;
  wire[2:0] CMeshDOR_3_io_outHeadFlit_priorityLevel;
  wire[2:0] CMeshDOR_3_io_result;
  wire[1:0] CMeshDOR_3_io_vcsAvailable_4;
  wire[1:0] CMeshDOR_3_io_vcsAvailable_3;
  wire[1:0] CMeshDOR_3_io_vcsAvailable_2;
  wire[1:0] CMeshDOR_3_io_vcsAvailable_1;
  wire[1:0] CMeshDOR_3_io_vcsAvailable_0;
  wire[2:0] VCRouterStateManagement_3_io_currentState;
  wire CreditGen_4_io_outCredit_grant;
  wire[54:0] RouterRegFile_4_io_readData;
  wire RouterRegFile_4_io_readValid;
  wire[54:0] RouterRegFile_4_io_readPipelineReg_1;
  wire[54:0] RouterRegFile_4_io_readPipelineReg_0;
  wire RouterRegFile_4_io_rvPipelineReg_1;
  wire RouterRegFile_4_io_rvPipelineReg_0;
  wire[15:0] CMeshDOR_4_io_outHeadFlit_packetID;
  wire CMeshDOR_4_io_outHeadFlit_isTail;
  wire CMeshDOR_4_io_outHeadFlit_vcPort;
  wire[3:0] CMeshDOR_4_io_outHeadFlit_packetType;
  wire[1:0] CMeshDOR_4_io_outHeadFlit_destination_2;
  wire[1:0] CMeshDOR_4_io_outHeadFlit_destination_1;
  wire[1:0] CMeshDOR_4_io_outHeadFlit_destination_0;
  wire[2:0] CMeshDOR_4_io_outHeadFlit_priorityLevel;
  wire[2:0] CMeshDOR_4_io_result;
  wire[1:0] CMeshDOR_4_io_vcsAvailable_4;
  wire[1:0] CMeshDOR_4_io_vcsAvailable_3;
  wire[1:0] CMeshDOR_4_io_vcsAvailable_2;
  wire[1:0] CMeshDOR_4_io_vcsAvailable_1;
  wire[1:0] CMeshDOR_4_io_vcsAvailable_0;
  wire[2:0] VCRouterStateManagement_4_io_currentState;
  wire CreditGen_5_io_outCredit_grant;
  wire[54:0] RouterRegFile_5_io_readData;
  wire RouterRegFile_5_io_readValid;
  wire[54:0] RouterRegFile_5_io_readPipelineReg_1;
  wire[54:0] RouterRegFile_5_io_readPipelineReg_0;
  wire RouterRegFile_5_io_rvPipelineReg_1;
  wire RouterRegFile_5_io_rvPipelineReg_0;
  wire[15:0] CMeshDOR_5_io_outHeadFlit_packetID;
  wire CMeshDOR_5_io_outHeadFlit_isTail;
  wire CMeshDOR_5_io_outHeadFlit_vcPort;
  wire[3:0] CMeshDOR_5_io_outHeadFlit_packetType;
  wire[1:0] CMeshDOR_5_io_outHeadFlit_destination_2;
  wire[1:0] CMeshDOR_5_io_outHeadFlit_destination_1;
  wire[1:0] CMeshDOR_5_io_outHeadFlit_destination_0;
  wire[2:0] CMeshDOR_5_io_outHeadFlit_priorityLevel;
  wire[2:0] CMeshDOR_5_io_result;
  wire[1:0] CMeshDOR_5_io_vcsAvailable_4;
  wire[1:0] CMeshDOR_5_io_vcsAvailable_3;
  wire[1:0] CMeshDOR_5_io_vcsAvailable_2;
  wire[1:0] CMeshDOR_5_io_vcsAvailable_1;
  wire[1:0] CMeshDOR_5_io_vcsAvailable_0;
  wire[2:0] VCRouterStateManagement_5_io_currentState;
  wire CreditGen_6_io_outCredit_grant;
  wire[54:0] RouterRegFile_6_io_readData;
  wire RouterRegFile_6_io_readValid;
  wire[54:0] RouterRegFile_6_io_readPipelineReg_1;
  wire[54:0] RouterRegFile_6_io_readPipelineReg_0;
  wire RouterRegFile_6_io_rvPipelineReg_1;
  wire RouterRegFile_6_io_rvPipelineReg_0;
  wire[15:0] CMeshDOR_6_io_outHeadFlit_packetID;
  wire CMeshDOR_6_io_outHeadFlit_isTail;
  wire CMeshDOR_6_io_outHeadFlit_vcPort;
  wire[3:0] CMeshDOR_6_io_outHeadFlit_packetType;
  wire[1:0] CMeshDOR_6_io_outHeadFlit_destination_2;
  wire[1:0] CMeshDOR_6_io_outHeadFlit_destination_1;
  wire[1:0] CMeshDOR_6_io_outHeadFlit_destination_0;
  wire[2:0] CMeshDOR_6_io_outHeadFlit_priorityLevel;
  wire[2:0] CMeshDOR_6_io_result;
  wire[1:0] CMeshDOR_6_io_vcsAvailable_4;
  wire[1:0] CMeshDOR_6_io_vcsAvailable_3;
  wire[1:0] CMeshDOR_6_io_vcsAvailable_2;
  wire[1:0] CMeshDOR_6_io_vcsAvailable_1;
  wire[1:0] CMeshDOR_6_io_vcsAvailable_0;
  wire[2:0] VCRouterStateManagement_6_io_currentState;
  wire CreditGen_7_io_outCredit_grant;
  wire[54:0] RouterRegFile_7_io_readData;
  wire RouterRegFile_7_io_readValid;
  wire[54:0] RouterRegFile_7_io_readPipelineReg_1;
  wire[54:0] RouterRegFile_7_io_readPipelineReg_0;
  wire RouterRegFile_7_io_rvPipelineReg_1;
  wire RouterRegFile_7_io_rvPipelineReg_0;
  wire[15:0] CMeshDOR_7_io_outHeadFlit_packetID;
  wire CMeshDOR_7_io_outHeadFlit_isTail;
  wire CMeshDOR_7_io_outHeadFlit_vcPort;
  wire[3:0] CMeshDOR_7_io_outHeadFlit_packetType;
  wire[1:0] CMeshDOR_7_io_outHeadFlit_destination_2;
  wire[1:0] CMeshDOR_7_io_outHeadFlit_destination_1;
  wire[1:0] CMeshDOR_7_io_outHeadFlit_destination_0;
  wire[2:0] CMeshDOR_7_io_outHeadFlit_priorityLevel;
  wire[2:0] CMeshDOR_7_io_result;
  wire[1:0] CMeshDOR_7_io_vcsAvailable_4;
  wire[1:0] CMeshDOR_7_io_vcsAvailable_3;
  wire[1:0] CMeshDOR_7_io_vcsAvailable_2;
  wire[1:0] CMeshDOR_7_io_vcsAvailable_1;
  wire[1:0] CMeshDOR_7_io_vcsAvailable_0;
  wire[2:0] VCRouterStateManagement_7_io_currentState;
  wire CreditGen_8_io_outCredit_grant;
  wire[54:0] RouterRegFile_8_io_readData;
  wire RouterRegFile_8_io_readValid;
  wire[54:0] RouterRegFile_8_io_readPipelineReg_1;
  wire[54:0] RouterRegFile_8_io_readPipelineReg_0;
  wire RouterRegFile_8_io_rvPipelineReg_1;
  wire RouterRegFile_8_io_rvPipelineReg_0;
  wire[15:0] CMeshDOR_8_io_outHeadFlit_packetID;
  wire CMeshDOR_8_io_outHeadFlit_isTail;
  wire CMeshDOR_8_io_outHeadFlit_vcPort;
  wire[3:0] CMeshDOR_8_io_outHeadFlit_packetType;
  wire[1:0] CMeshDOR_8_io_outHeadFlit_destination_2;
  wire[1:0] CMeshDOR_8_io_outHeadFlit_destination_1;
  wire[1:0] CMeshDOR_8_io_outHeadFlit_destination_0;
  wire[2:0] CMeshDOR_8_io_outHeadFlit_priorityLevel;
  wire[2:0] CMeshDOR_8_io_result;
  wire[1:0] CMeshDOR_8_io_vcsAvailable_4;
  wire[1:0] CMeshDOR_8_io_vcsAvailable_3;
  wire[1:0] CMeshDOR_8_io_vcsAvailable_2;
  wire[1:0] CMeshDOR_8_io_vcsAvailable_1;
  wire[1:0] CMeshDOR_8_io_vcsAvailable_0;
  wire[2:0] VCRouterStateManagement_8_io_currentState;
  wire CreditGen_9_io_outCredit_grant;
  wire[54:0] RouterRegFile_9_io_readData;
  wire RouterRegFile_9_io_readValid;
  wire[54:0] RouterRegFile_9_io_readPipelineReg_1;
  wire[54:0] RouterRegFile_9_io_readPipelineReg_0;
  wire RouterRegFile_9_io_rvPipelineReg_1;
  wire RouterRegFile_9_io_rvPipelineReg_0;
  wire[15:0] CMeshDOR_9_io_outHeadFlit_packetID;
  wire CMeshDOR_9_io_outHeadFlit_isTail;
  wire CMeshDOR_9_io_outHeadFlit_vcPort;
  wire[3:0] CMeshDOR_9_io_outHeadFlit_packetType;
  wire[1:0] CMeshDOR_9_io_outHeadFlit_destination_2;
  wire[1:0] CMeshDOR_9_io_outHeadFlit_destination_1;
  wire[1:0] CMeshDOR_9_io_outHeadFlit_destination_0;
  wire[2:0] CMeshDOR_9_io_outHeadFlit_priorityLevel;
  wire[2:0] CMeshDOR_9_io_result;
  wire[1:0] CMeshDOR_9_io_vcsAvailable_4;
  wire[1:0] CMeshDOR_9_io_vcsAvailable_3;
  wire[1:0] CMeshDOR_9_io_vcsAvailable_2;
  wire[1:0] CMeshDOR_9_io_vcsAvailable_1;
  wire[1:0] CMeshDOR_9_io_vcsAvailable_0;
  wire[2:0] VCRouterStateManagement_9_io_currentState;
  wire CreditCon_io_outCredit;
  wire CreditCon_1_io_outCredit;
  wire CreditCon_2_io_outCredit;
  wire CreditCon_3_io_outCredit;
  wire CreditCon_4_io_outCredit;
  wire CreditCon_5_io_outCredit;
  wire CreditCon_6_io_outCredit;
  wire CreditCon_7_io_outCredit;
  wire CreditCon_8_io_outCredit;
  wire CreditCon_9_io_outCredit;
  wire[54:0] switch_io_outPorts_4_x;
  wire[54:0] switch_io_outPorts_3_x;
  wire[54:0] switch_io_outPorts_2_x;
  wire[54:0] switch_io_outPorts_1_x;
  wire[54:0] switch_io_outPorts_0_x;
  wire swAllocator_io_requests_4_9_grant;
  wire swAllocator_io_requests_4_8_grant;
  wire swAllocator_io_requests_4_7_grant;
  wire swAllocator_io_requests_4_6_grant;
  wire swAllocator_io_requests_4_5_grant;
  wire swAllocator_io_requests_4_4_grant;
  wire swAllocator_io_requests_4_3_grant;
  wire swAllocator_io_requests_4_2_grant;
  wire swAllocator_io_requests_4_1_grant;
  wire swAllocator_io_requests_4_0_grant;
  wire swAllocator_io_requests_3_9_grant;
  wire swAllocator_io_requests_3_8_grant;
  wire swAllocator_io_requests_3_7_grant;
  wire swAllocator_io_requests_3_6_grant;
  wire swAllocator_io_requests_3_5_grant;
  wire swAllocator_io_requests_3_4_grant;
  wire swAllocator_io_requests_3_3_grant;
  wire swAllocator_io_requests_3_2_grant;
  wire swAllocator_io_requests_3_1_grant;
  wire swAllocator_io_requests_3_0_grant;
  wire swAllocator_io_requests_2_9_grant;
  wire swAllocator_io_requests_2_8_grant;
  wire swAllocator_io_requests_2_7_grant;
  wire swAllocator_io_requests_2_6_grant;
  wire swAllocator_io_requests_2_5_grant;
  wire swAllocator_io_requests_2_4_grant;
  wire swAllocator_io_requests_2_3_grant;
  wire swAllocator_io_requests_2_2_grant;
  wire swAllocator_io_requests_2_1_grant;
  wire swAllocator_io_requests_2_0_grant;
  wire swAllocator_io_requests_1_9_grant;
  wire swAllocator_io_requests_1_8_grant;
  wire swAllocator_io_requests_1_7_grant;
  wire swAllocator_io_requests_1_6_grant;
  wire swAllocator_io_requests_1_5_grant;
  wire swAllocator_io_requests_1_4_grant;
  wire swAllocator_io_requests_1_3_grant;
  wire swAllocator_io_requests_1_2_grant;
  wire swAllocator_io_requests_1_1_grant;
  wire swAllocator_io_requests_1_0_grant;
  wire swAllocator_io_requests_0_9_grant;
  wire swAllocator_io_requests_0_8_grant;
  wire swAllocator_io_requests_0_7_grant;
  wire swAllocator_io_requests_0_6_grant;
  wire swAllocator_io_requests_0_5_grant;
  wire swAllocator_io_requests_0_4_grant;
  wire swAllocator_io_requests_0_3_grant;
  wire swAllocator_io_requests_0_2_grant;
  wire swAllocator_io_requests_0_1_grant;
  wire swAllocator_io_requests_0_0_grant;
  wire[3:0] swAllocator_io_chosens_4;
  wire[3:0] swAllocator_io_chosens_3;
  wire[3:0] swAllocator_io_chosens_2;
  wire[3:0] swAllocator_io_chosens_1;
  wire[3:0] swAllocator_io_chosens_0;
  wire vcAllocator_io_resources_9_valid;
  wire vcAllocator_io_resources_8_valid;
  wire vcAllocator_io_resources_7_valid;
  wire vcAllocator_io_resources_6_valid;
  wire vcAllocator_io_resources_5_valid;
  wire vcAllocator_io_resources_4_valid;
  wire vcAllocator_io_resources_3_valid;
  wire vcAllocator_io_resources_2_valid;
  wire vcAllocator_io_resources_1_valid;
  wire vcAllocator_io_resources_0_valid;
  wire[3:0] vcAllocator_io_chosens_9;
  wire[3:0] vcAllocator_io_chosens_8;
  wire[3:0] vcAllocator_io_chosens_7;
  wire[3:0] vcAllocator_io_chosens_6;
  wire[3:0] vcAllocator_io_chosens_5;
  wire[3:0] vcAllocator_io_chosens_4;
  wire[3:0] vcAllocator_io_chosens_3;
  wire[3:0] vcAllocator_io_chosens_2;
  wire[3:0] vcAllocator_io_chosens_1;
  wire[3:0] vcAllocator_io_chosens_0;
  wire RouterBuffer_io_enq_ready;
  wire RouterBuffer_io_deq_valid;
  wire[54:0] RouterBuffer_io_deq_bits_x;
  wire[54:0] ReplaceVCPort_io_newFlit_x;
  wire RouterBuffer_1_io_enq_ready;
  wire RouterBuffer_1_io_deq_valid;
  wire[54:0] RouterBuffer_1_io_deq_bits_x;
  wire[54:0] ReplaceVCPort_1_io_newFlit_x;
  wire RouterBuffer_2_io_enq_ready;
  wire RouterBuffer_2_io_deq_valid;
  wire[54:0] RouterBuffer_2_io_deq_bits_x;
  wire[54:0] ReplaceVCPort_2_io_newFlit_x;
  wire RouterBuffer_3_io_enq_ready;
  wire RouterBuffer_3_io_deq_valid;
  wire[54:0] RouterBuffer_3_io_deq_bits_x;
  wire[54:0] ReplaceVCPort_3_io_newFlit_x;
  wire RouterBuffer_4_io_enq_ready;
  wire RouterBuffer_4_io_deq_valid;
  wire[54:0] RouterBuffer_4_io_deq_bits_x;
  wire[54:0] ReplaceVCPort_4_io_newFlit_x;
  wire RouterBuffer_5_io_enq_ready;
  wire RouterBuffer_5_io_deq_valid;
  wire[54:0] RouterBuffer_5_io_deq_bits_x;
  wire[54:0] ReplaceVCPort_5_io_newFlit_x;
  wire RouterBuffer_6_io_enq_ready;
  wire RouterBuffer_6_io_deq_valid;
  wire[54:0] RouterBuffer_6_io_deq_bits_x;
  wire[54:0] ReplaceVCPort_6_io_newFlit_x;
  wire RouterBuffer_7_io_enq_ready;
  wire RouterBuffer_7_io_deq_valid;
  wire[54:0] RouterBuffer_7_io_deq_bits_x;
  wire[54:0] ReplaceVCPort_7_io_newFlit_x;
  wire RouterBuffer_8_io_enq_ready;
  wire RouterBuffer_8_io_deq_valid;
  wire[54:0] RouterBuffer_8_io_deq_bits_x;
  wire[54:0] ReplaceVCPort_8_io_newFlit_x;
  wire RouterBuffer_9_io_enq_ready;
  wire RouterBuffer_9_io_deq_valid;
  wire[54:0] RouterBuffer_9_io_deq_bits_x;
  wire[54:0] ReplaceVCPort_9_io_newFlit_x;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    T0 = 1'b0;
    T17 = 1'b0;
    T22 = 1'b0;
    T39 = 1'b0;
    T44 = 1'b0;
    T61 = 1'b0;
    T66 = 1'b0;
    T83 = 1'b0;
    T88 = 1'b0;
    T105 = 1'b0;
    T110 = 1'b0;
    T127 = 1'b0;
    T132 = 1'b0;
    T149 = 1'b0;
    T154 = 1'b0;
    T171 = 1'b0;
    T176 = 1'b0;
    T193 = 1'b0;
    T198 = 1'b0;
    T215 = 1'b0;
    R282 = {2{1'b0}};
    R295 = {1{1'b0}};
    R349 = {1{1'b0}};
    R426 = {2{1'b0}};
    R439 = {1{1'b0}};
    R493 = {1{1'b0}};
    R570 = {2{1'b0}};
    R583 = {1{1'b0}};
    R637 = {1{1'b0}};
    R714 = {2{1'b0}};
    R727 = {1{1'b0}};
    R781 = {1{1'b0}};
    R858 = {2{1'b0}};
    R871 = {1{1'b0}};
    R925 = {1{1'b0}};
    R1002 = {2{1'b0}};
    R1015 = {1{1'b0}};
    R1069 = {1{1'b0}};
    R1146 = {2{1'b0}};
    R1159 = {1{1'b0}};
    R1213 = {1{1'b0}};
    R1290 = {2{1'b0}};
    R1303 = {1{1'b0}};
    R1357 = {1{1'b0}};
    R1434 = {2{1'b0}};
    R1447 = {1{1'b0}};
    R1501 = {1{1'b0}};
    R1578 = {2{1'b0}};
    R1591 = {1{1'b0}};
    R1645 = {1{1'b0}};
    validVCs_0_0 = {1{1'b0}};
    R2176 = {1{1'b0}};
    R2181 = {1{1'b0}};
    validVCs_0_1 = {1{1'b0}};
    R2186 = {1{1'b0}};
    R2191 = {1{1'b0}};
    validVCs_0_2 = {1{1'b0}};
    R2196 = {1{1'b0}};
    R2201 = {1{1'b0}};
    validVCs_0_3 = {1{1'b0}};
    R2206 = {1{1'b0}};
    R2211 = {1{1'b0}};
    validVCs_0_4 = {1{1'b0}};
    R2216 = {1{1'b0}};
    R2221 = {1{1'b0}};
    validVCs_1_0 = {1{1'b0}};
    R2226 = {1{1'b0}};
    R2231 = {1{1'b0}};
    validVCs_1_1 = {1{1'b0}};
    R2236 = {1{1'b0}};
    R2241 = {1{1'b0}};
    validVCs_1_2 = {1{1'b0}};
    R2246 = {1{1'b0}};
    R2251 = {1{1'b0}};
    validVCs_1_3 = {1{1'b0}};
    R2256 = {1{1'b0}};
    R2261 = {1{1'b0}};
    validVCs_1_4 = {1{1'b0}};
    R2266 = {1{1'b0}};
    R2271 = {1{1'b0}};
    validVCs_2_0 = {1{1'b0}};
    R2276 = {1{1'b0}};
    R2281 = {1{1'b0}};
    validVCs_2_1 = {1{1'b0}};
    R2286 = {1{1'b0}};
    R2291 = {1{1'b0}};
    validVCs_2_2 = {1{1'b0}};
    R2296 = {1{1'b0}};
    R2301 = {1{1'b0}};
    validVCs_2_3 = {1{1'b0}};
    R2306 = {1{1'b0}};
    R2311 = {1{1'b0}};
    validVCs_2_4 = {1{1'b0}};
    R2316 = {1{1'b0}};
    R2321 = {1{1'b0}};
    validVCs_3_0 = {1{1'b0}};
    R2326 = {1{1'b0}};
    R2331 = {1{1'b0}};
    validVCs_3_1 = {1{1'b0}};
    R2336 = {1{1'b0}};
    R2341 = {1{1'b0}};
    validVCs_3_2 = {1{1'b0}};
    R2346 = {1{1'b0}};
    R2351 = {1{1'b0}};
    validVCs_3_3 = {1{1'b0}};
    R2356 = {1{1'b0}};
    R2361 = {1{1'b0}};
    validVCs_3_4 = {1{1'b0}};
    R2366 = {1{1'b0}};
    R2371 = {1{1'b0}};
    validVCs_4_0 = {1{1'b0}};
    R2376 = {1{1'b0}};
    R2381 = {1{1'b0}};
    validVCs_4_1 = {1{1'b0}};
    R2386 = {1{1'b0}};
    R2391 = {1{1'b0}};
    validVCs_4_2 = {1{1'b0}};
    R2396 = {1{1'b0}};
    R2401 = {1{1'b0}};
    validVCs_4_3 = {1{1'b0}};
    R2406 = {1{1'b0}};
    R2411 = {1{1'b0}};
    validVCs_4_4 = {1{1'b0}};
    R2416 = {1{1'b0}};
    R2421 = {1{1'b0}};
    validVCs_5_0 = {1{1'b0}};
    R2426 = {1{1'b0}};
    R2431 = {1{1'b0}};
    validVCs_5_1 = {1{1'b0}};
    R2436 = {1{1'b0}};
    R2441 = {1{1'b0}};
    validVCs_5_2 = {1{1'b0}};
    R2446 = {1{1'b0}};
    R2451 = {1{1'b0}};
    validVCs_5_3 = {1{1'b0}};
    R2456 = {1{1'b0}};
    R2461 = {1{1'b0}};
    validVCs_5_4 = {1{1'b0}};
    R2466 = {1{1'b0}};
    R2471 = {1{1'b0}};
    validVCs_6_0 = {1{1'b0}};
    R2476 = {1{1'b0}};
    R2481 = {1{1'b0}};
    validVCs_6_1 = {1{1'b0}};
    R2486 = {1{1'b0}};
    R2491 = {1{1'b0}};
    validVCs_6_2 = {1{1'b0}};
    R2496 = {1{1'b0}};
    R2501 = {1{1'b0}};
    validVCs_6_3 = {1{1'b0}};
    R2506 = {1{1'b0}};
    R2511 = {1{1'b0}};
    validVCs_6_4 = {1{1'b0}};
    R2516 = {1{1'b0}};
    R2521 = {1{1'b0}};
    validVCs_7_0 = {1{1'b0}};
    R2526 = {1{1'b0}};
    R2531 = {1{1'b0}};
    validVCs_7_1 = {1{1'b0}};
    R2536 = {1{1'b0}};
    R2541 = {1{1'b0}};
    validVCs_7_2 = {1{1'b0}};
    R2546 = {1{1'b0}};
    R2551 = {1{1'b0}};
    validVCs_7_3 = {1{1'b0}};
    R2556 = {1{1'b0}};
    R2561 = {1{1'b0}};
    validVCs_7_4 = {1{1'b0}};
    R2566 = {1{1'b0}};
    R2571 = {1{1'b0}};
    validVCs_8_0 = {1{1'b0}};
    R2576 = {1{1'b0}};
    R2581 = {1{1'b0}};
    validVCs_8_1 = {1{1'b0}};
    R2586 = {1{1'b0}};
    R2591 = {1{1'b0}};
    validVCs_8_2 = {1{1'b0}};
    R2596 = {1{1'b0}};
    R2601 = {1{1'b0}};
    validVCs_8_3 = {1{1'b0}};
    R2606 = {1{1'b0}};
    R2611 = {1{1'b0}};
    validVCs_8_4 = {1{1'b0}};
    R2616 = {1{1'b0}};
    R2621 = {1{1'b0}};
    validVCs_9_0 = {1{1'b0}};
    R2626 = {1{1'b0}};
    R2631 = {1{1'b0}};
    validVCs_9_1 = {1{1'b0}};
    R2636 = {1{1'b0}};
    R2641 = {1{1'b0}};
    validVCs_9_2 = {1{1'b0}};
    R2646 = {1{1'b0}};
    R2651 = {1{1'b0}};
    validVCs_9_3 = {1{1'b0}};
    R2656 = {1{1'b0}};
    R2661 = {1{1'b0}};
    validVCs_9_4 = {1{1'b0}};
    R2666 = {1{1'b0}};
    R2671 = {1{1'b0}};
    R2675 = {1{1'b0}};
    R2683 = {1{1'b0}};
    R2688 = {1{1'b0}};
    R2689 = {1{1'b0}};
    R2697 = {1{1'b0}};
    R2702 = {1{1'b0}};
    R2703 = {1{1'b0}};
    R2711 = {1{1'b0}};
    R2716 = {1{1'b0}};
    R2717 = {1{1'b0}};
    R2725 = {1{1'b0}};
    R2730 = {1{1'b0}};
    R2731 = {1{1'b0}};
    R2739 = {1{1'b0}};
    R2744 = {1{1'b0}};
    R2745 = {1{1'b0}};
    R2753 = {1{1'b0}};
    R2758 = {1{1'b0}};
    R2759 = {1{1'b0}};
    R2767 = {1{1'b0}};
    R2772 = {1{1'b0}};
    R2773 = {1{1'b0}};
    R2781 = {1{1'b0}};
    R2786 = {1{1'b0}};
    R2787 = {1{1'b0}};
    R2795 = {1{1'b0}};
    R2800 = {1{1'b0}};
    R2801 = {1{1'b0}};
    R2809 = {1{1'b0}};
    R2814 = {1{1'b0}};
    R3097 = {1{1'b0}};
    R3098 = {2{1'b0}};
    R3100 = {1{1'b0}};
    R3101 = {2{1'b0}};
    R3103 = {1{1'b0}};
    R3104 = {2{1'b0}};
    R3106 = {1{1'b0}};
    R3107 = {2{1'b0}};
    R3109 = {1{1'b0}};
    R3110 = {2{1'b0}};
  end
// synthesis translate_on
`endif

`ifndef SYNTHESIS
// synthesis translate_off
//  assign io_counters_0_counterIndex = {1{1'b0}};
//  assign io_counters_1_counterIndex = {1{1'b0}};
//  assign io_counters_1_counterVal = {1{1'b0}};
// synthesis translate_on
`endif
  assign T1 = T2 | reset;
  assign T2 = T13 | T3;
  assign T3 = ~ T4;
  assign T4 = T5 == 1'h1;
  assign T5 = T6;
  assign T6 = T11 ? T9 : T7;
  assign T7 = T8[6'h24:6'h24];
  assign T8 = io_inChannels_4_flit_x[6'h36:1'h1];
  assign T9 = T10[4'hd:4'hd];
  assign T10 = io_inChannels_4_flit_x[5'h1f:1'h1];
  assign T11 = T12 == 1'h1;
  assign T12 = io_inChannels_4_flit_x[1'h0:1'h0];
  assign T13 = T15 | T14;
  assign T14 = ~ io_inChannels_4_flitValid;
  assign T15 = T16 & T4;
  assign T16 = RouterBuffer_9_io_enq_ready & io_inChannels_4_flitValid;
  assign T18 = T19 | reset;
  assign T19 = T21 | T20;
  assign T20 = T379 & T4;
  assign T21 = ~ T379;
  assign T23 = T24 | reset;
  assign T24 = T35 | T25;
  assign T25 = ~ T26;
  assign T26 = T27 == 1'h0;
  assign T27 = T28;
  assign T28 = T33 ? T31 : T29;
  assign T29 = T30[6'h24:6'h24];
  assign T30 = io_inChannels_4_flit_x[6'h36:1'h1];
  assign T31 = T32[4'hd:4'hd];
  assign T32 = io_inChannels_4_flit_x[5'h1f:1'h1];
  assign T33 = T34 == 1'h1;
  assign T34 = io_inChannels_4_flit_x[1'h0:1'h0];
  assign T35 = T37 | T36;
  assign T36 = ~ io_inChannels_4_flitValid;
  assign T37 = T38 & T26;
  assign T38 = RouterBuffer_8_io_enq_ready & io_inChannels_4_flitValid;
  assign T40 = T41 | reset;
  assign T41 = T43 | T42;
  assign T42 = T523 & T26;
  assign T43 = ~ T523;
  assign T45 = T46 | reset;
  assign T46 = T57 | T47;
  assign T47 = ~ T48;
  assign T48 = T49 == 1'h1;
  assign T49 = T50;
  assign T50 = T55 ? T53 : T51;
  assign T51 = T52[6'h24:6'h24];
  assign T52 = io_inChannels_3_flit_x[6'h36:1'h1];
  assign T53 = T54[4'hd:4'hd];
  assign T54 = io_inChannels_3_flit_x[5'h1f:1'h1];
  assign T55 = T56 == 1'h1;
  assign T56 = io_inChannels_3_flit_x[1'h0:1'h0];
  assign T57 = T59 | T58;
  assign T58 = ~ io_inChannels_3_flitValid;
  assign T59 = T60 & T48;
  assign T60 = RouterBuffer_7_io_enq_ready & io_inChannels_3_flitValid;
  assign T62 = T63 | reset;
  assign T63 = T65 | T64;
  assign T64 = T667 & T48;
  assign T65 = ~ T667;
  assign T67 = T68 | reset;
  assign T68 = T79 | T69;
  assign T69 = ~ T70;
  assign T70 = T71 == 1'h0;
  assign T71 = T72;
  assign T72 = T77 ? T75 : T73;
  assign T73 = T74[6'h24:6'h24];
  assign T74 = io_inChannels_3_flit_x[6'h36:1'h1];
  assign T75 = T76[4'hd:4'hd];
  assign T76 = io_inChannels_3_flit_x[5'h1f:1'h1];
  assign T77 = T78 == 1'h1;
  assign T78 = io_inChannels_3_flit_x[1'h0:1'h0];
  assign T79 = T81 | T80;
  assign T80 = ~ io_inChannels_3_flitValid;
  assign T81 = T82 & T70;
  assign T82 = RouterBuffer_6_io_enq_ready & io_inChannels_3_flitValid;
  assign T84 = T85 | reset;
  assign T85 = T87 | T86;
  assign T86 = T811 & T70;
  assign T87 = ~ T811;
  assign T89 = T90 | reset;
  assign T90 = T101 | T91;
  assign T91 = ~ T92;
  assign T92 = T93 == 1'h1;
  assign T93 = T94;
  assign T94 = T99 ? T97 : T95;
  assign T95 = T96[6'h24:6'h24];
  assign T96 = io_inChannels_2_flit_x[6'h36:1'h1];
  assign T97 = T98[4'hd:4'hd];
  assign T98 = io_inChannels_2_flit_x[5'h1f:1'h1];
  assign T99 = T100 == 1'h1;
  assign T100 = io_inChannels_2_flit_x[1'h0:1'h0];
  assign T101 = T103 | T102;
  assign T102 = ~ io_inChannels_2_flitValid;
  assign T103 = T104 & T92;
  assign T104 = RouterBuffer_5_io_enq_ready & io_inChannels_2_flitValid;
  assign T106 = T107 | reset;
  assign T107 = T109 | T108;
  assign T108 = T955 & T92;
  assign T109 = ~ T955;
  assign T111 = T112 | reset;
  assign T112 = T123 | T113;
  assign T113 = ~ T114;
  assign T114 = T115 == 1'h0;
  assign T115 = T116;
  assign T116 = T121 ? T119 : T117;
  assign T117 = T118[6'h24:6'h24];
  assign T118 = io_inChannels_2_flit_x[6'h36:1'h1];
  assign T119 = T120[4'hd:4'hd];
  assign T120 = io_inChannels_2_flit_x[5'h1f:1'h1];
  assign T121 = T122 == 1'h1;
  assign T122 = io_inChannels_2_flit_x[1'h0:1'h0];
  assign T123 = T125 | T124;
  assign T124 = ~ io_inChannels_2_flitValid;
  assign T125 = T126 & T114;
  assign T126 = RouterBuffer_4_io_enq_ready & io_inChannels_2_flitValid;
  assign T128 = T129 | reset;
  assign T129 = T131 | T130;
  assign T130 = T1099 & T114;
  assign T131 = ~ T1099;
  assign T133 = T134 | reset;
  assign T134 = T145 | T135;
  assign T135 = ~ T136;
  assign T136 = T137 == 1'h1;
  assign T137 = T138;
  assign T138 = T143 ? T141 : T139;
  assign T139 = T140[6'h24:6'h24];
  assign T140 = io_inChannels_1_flit_x[6'h36:1'h1];
  assign T141 = T142[4'hd:4'hd];
  assign T142 = io_inChannels_1_flit_x[5'h1f:1'h1];
  assign T143 = T144 == 1'h1;
  assign T144 = io_inChannels_1_flit_x[1'h0:1'h0];
  assign T145 = T147 | T146;
  assign T146 = ~ io_inChannels_1_flitValid;
  assign T147 = T148 & T136;
  assign T148 = RouterBuffer_3_io_enq_ready & io_inChannels_1_flitValid;
  assign T150 = T151 | reset;
  assign T151 = T153 | T152;
  assign T152 = T1243 & T136;
  assign T153 = ~ T1243;
  assign T155 = T156 | reset;
  assign T156 = T167 | T157;
  assign T157 = ~ T158;
  assign T158 = T159 == 1'h0;
  assign T159 = T160;
  assign T160 = T165 ? T163 : T161;
  assign T161 = T162[6'h24:6'h24];
  assign T162 = io_inChannels_1_flit_x[6'h36:1'h1];
  assign T163 = T164[4'hd:4'hd];
  assign T164 = io_inChannels_1_flit_x[5'h1f:1'h1];
  assign T165 = T166 == 1'h1;
  assign T166 = io_inChannels_1_flit_x[1'h0:1'h0];
  assign T167 = T169 | T168;
  assign T168 = ~ io_inChannels_1_flitValid;
  assign T169 = T170 & T158;
  assign T170 = RouterBuffer_2_io_enq_ready & io_inChannels_1_flitValid;
  assign T172 = T173 | reset;
  assign T173 = T175 | T174;
  assign T174 = T1387 & T158;
  assign T175 = ~ T1387;
  assign T177 = T178 | reset;
  assign T178 = T189 | T179;
  assign T179 = ~ T180;
  assign T180 = T181 == 1'h1;
  assign T181 = T182;
  assign T182 = T187 ? T185 : T183;
  assign T183 = T184[6'h24:6'h24];
  assign T184 = io_inChannels_0_flit_x[6'h36:1'h1];
  assign T185 = T186[4'hd:4'hd];
  assign T186 = io_inChannels_0_flit_x[5'h1f:1'h1];
  assign T187 = T188 == 1'h1;
  assign T188 = io_inChannels_0_flit_x[1'h0:1'h0];
  assign T189 = T191 | T190;
  assign T190 = ~ io_inChannels_0_flitValid;
  assign T191 = T192 & T180;
  assign T192 = RouterBuffer_1_io_enq_ready & io_inChannels_0_flitValid;
  assign T194 = T195 | reset;
  assign T195 = T197 | T196;
  assign T196 = T1531 & T180;
  assign T197 = ~ T1531;
  assign T199 = T200 | reset;
  assign T200 = T211 | T201;
  assign T201 = ~ T202;
  assign T202 = T203 == 1'h0;
  assign T203 = T204;
  assign T204 = T209 ? T207 : T205;
  assign T205 = T206[6'h24:6'h24];
  assign T206 = io_inChannels_0_flit_x[6'h36:1'h1];
  assign T207 = T208[4'hd:4'hd];
  assign T208 = io_inChannels_0_flit_x[5'h1f:1'h1];
  assign T209 = T210 == 1'h1;
  assign T210 = io_inChannels_0_flit_x[1'h0:1'h0];
  assign T211 = T213 | T212;
  assign T212 = ~ io_inChannels_0_flitValid;
  assign T213 = T214 & T202;
  assign T214 = RouterBuffer_io_enq_ready & io_inChannels_0_flitValid;
  assign T216 = T217 | reset;
  assign T217 = T219 | T218;
  assign T218 = T1675 & T202;
  assign T219 = ~ T1675;
  assign T220 = T1722 & T221;
  assign T221 = T222 == 1'h1;
  assign T222 = T223;
  assign T223 = T228 ? T226 : T224;
  assign T224 = T225[6'h24:6'h24];
  assign T225 = switch_io_outPorts_4_x[6'h36:1'h1];
  assign T226 = T227[4'hd:4'hd];
  assign T227 = switch_io_outPorts_4_x[5'h1f:1'h1];
  assign T228 = T229 == 1'h1;
  assign T229 = switch_io_outPorts_4_x[1'h0:1'h0];
  assign T230 = T1722 & T231;
  assign T231 = T222 == 1'h0;
  assign T232 = T1905 & T233;
  assign T233 = T234 == 1'h1;
  assign T234 = T235;
  assign T235 = T240 ? T238 : T236;
  assign T236 = T237[6'h24:6'h24];
  assign T237 = switch_io_outPorts_3_x[6'h36:1'h1];
  assign T238 = T239[4'hd:4'hd];
  assign T239 = switch_io_outPorts_3_x[5'h1f:1'h1];
  assign T240 = T241 == 1'h1;
  assign T241 = switch_io_outPorts_3_x[1'h0:1'h0];
  assign T242 = T1905 & T243;
  assign T243 = T234 == 1'h0;
  assign T244 = T1968 & T245;
  assign T245 = T246 == 1'h1;
  assign T246 = T247;
  assign T247 = T252 ? T250 : T248;
  assign T248 = T249[6'h24:6'h24];
  assign T249 = switch_io_outPorts_2_x[6'h36:1'h1];
  assign T250 = T251[4'hd:4'hd];
  assign T251 = switch_io_outPorts_2_x[5'h1f:1'h1];
  assign T252 = T253 == 1'h1;
  assign T253 = switch_io_outPorts_2_x[1'h0:1'h0];
  assign T254 = T1968 & T255;
  assign T255 = T246 == 1'h0;
  assign T256 = T2031 & T257;
  assign T257 = T258 == 1'h1;
  assign T258 = T259;
  assign T259 = T264 ? T262 : T260;
  assign T260 = T261[6'h24:6'h24];
  assign T261 = switch_io_outPorts_1_x[6'h36:1'h1];
  assign T262 = T263[4'hd:4'hd];
  assign T263 = switch_io_outPorts_1_x[5'h1f:1'h1];
  assign T264 = T265 == 1'h1;
  assign T265 = switch_io_outPorts_1_x[1'h0:1'h0];
  assign T266 = T2031 & T267;
  assign T267 = T258 == 1'h0;
  assign T268 = T2094 & T269;
  assign T269 = T270 == 1'h1;
  assign T270 = T271;
  assign T271 = T276 ? T274 : T272;
  assign T272 = T273[6'h24:6'h24];
  assign T273 = switch_io_outPorts_0_x[6'h36:1'h1];
  assign T274 = T275[4'hd:4'hd];
  assign T275 = switch_io_outPorts_0_x[5'h1f:1'h1];
  assign T276 = T277 == 1'h1;
  assign T277 = switch_io_outPorts_0_x[1'h0:1'h0];
  assign T278 = T2094 & T279;
  assign T279 = T270 == 1'h0;
  assign T280 = T281;
  assign T281 = io_inChannels_4_flit_x;
  assign T3112 = R282[1'h0:1'h0];
  assign T3113 = reset ? 55'h0 : T283;
  assign T283 = T284 ? T3114 : R282;
  assign T3114 = {51'h0, vcAllocator_io_chosens_9};
  assign T284 = T285 & vcAllocator_io_resources_9_valid;
  assign T285 = VCRouterStateManagement_9_io_currentState == 3'h2;
  assign T286 = T287;
  assign T287 = RouterBuffer_9_io_deq_bits_x;
  assign T288 = T300 | T289;
  assign T289 = T290 == 2'h1;
  assign T290 = T299 ? VCRouterOutputStateManagement_4_io_currentState : T291;
  assign T291 = T298 ? T296 : T292;
  assign T292 = T293 ? VCRouterOutputStateManagement_1_io_currentState : VCRouterOutputStateManagement_io_currentState;
  assign T293 = T294[1'h0:1'h0];
  assign T294 = R295;
  assign T3115 = reset ? 3'h0 : CMeshDOR_9_io_result;
  assign T296 = T297 ? VCRouterOutputStateManagement_3_io_currentState : VCRouterOutputStateManagement_2_io_currentState;
  assign T297 = T294[1'h0:1'h0];
  assign T298 = T294[1'h1:1'h1];
  assign T299 = T294[2'h2:2'h2];
  assign T300 = T290 == 2'h2;
  assign T301 = T319 ? T311 : T302;
  assign T302 = T310 ? creditConsReady_4_0 : T303;
  assign T303 = T309 ? T307 : T304;
  assign T304 = T305 ? creditConsReady_1_0 : creditConsReady_0_0;
  assign creditConsReady_0_0 = CreditCon_io_outCredit;
  assign creditConsReady_1_0 = CreditCon_2_io_outCredit;
  assign T305 = T306[1'h0:1'h0];
  assign T306 = R295;
  assign T307 = T308 ? creditConsReady_3_0 : creditConsReady_2_0;
  assign creditConsReady_2_0 = CreditCon_4_io_outCredit;
  assign creditConsReady_3_0 = CreditCon_6_io_outCredit;
  assign T308 = T306[1'h0:1'h0];
  assign T309 = T306[1'h1:1'h1];
  assign creditConsReady_4_0 = CreditCon_8_io_outCredit;
  assign T310 = T306[2'h2:2'h2];
  assign T311 = T318 ? creditConsReady_4_1 : T312;
  assign T312 = T317 ? T315 : T313;
  assign T313 = T314 ? creditConsReady_1_1 : creditConsReady_0_1;
  assign creditConsReady_0_1 = CreditCon_1_io_outCredit;
  assign creditConsReady_1_1 = CreditCon_3_io_outCredit;
  assign T314 = T306[1'h0:1'h0];
  assign T315 = T316 ? creditConsReady_3_1 : creditConsReady_2_1;
  assign creditConsReady_2_1 = CreditCon_5_io_outCredit;
  assign creditConsReady_3_1 = CreditCon_7_io_outCredit;
  assign T316 = T306[1'h0:1'h0];
  assign T317 = T306[1'h1:1'h1];
  assign creditConsReady_4_1 = CreditCon_9_io_outCredit;
  assign T318 = T306[2'h2:2'h2];
  assign T319 = T3116;
  assign T3116 = R282[1'h0:1'h0];
  assign T320 = T331 & T321;
  assign T321 = T322 == 4'h9;
  assign T322 = T330 ? swAllocator_io_chosens_4 : T323;
  assign T323 = T329 ? T327 : T324;
  assign T324 = T325 ? swAllocator_io_chosens_1 : swAllocator_io_chosens_0;
  assign T325 = T326[1'h0:1'h0];
  assign T326 = R295;
  assign T327 = T328 ? swAllocator_io_chosens_3 : swAllocator_io_chosens_2;
  assign T328 = T326[1'h0:1'h0];
  assign T329 = T326[1'h1:1'h1];
  assign T330 = T326[2'h2:2'h2];
  assign T331 = T339 ? swAllocator_io_requests_4_9_grant : T332;
  assign T332 = T338 ? T336 : T333;
  assign T333 = T334 ? swAllocator_io_requests_1_9_grant : swAllocator_io_requests_0_9_grant;
  assign T334 = T335[1'h0:1'h0];
  assign T335 = R295;
  assign T336 = T337 ? swAllocator_io_requests_3_9_grant : swAllocator_io_requests_2_9_grant;
  assign T337 = T335[1'h0:1'h0];
  assign T338 = T335[1'h1:1'h1];
  assign T339 = T335[2'h2:2'h2];
  assign T340 = RouterBuffer_9_io_deq_valid & T341;
  assign T341 = T342;
  assign T342 = T347 ? T345 : T343;
  assign T343 = T344[6'h25:6'h25];
  assign T344 = RouterBuffer_9_io_deq_bits_x[6'h36:1'h1];
  assign T345 = T346[4'he:4'he];
  assign T346 = RouterBuffer_9_io_deq_bits_x[5'h1f:1'h1];
  assign T347 = T348 == 1'h1;
  assign T348 = RouterBuffer_9_io_deq_bits_x[1'h0:1'h0];
  assign T3117 = reset ? 1'h0 : RouterBuffer_9_io_deq_valid;
  assign T350 = T351[2'h2:1'h0];
  assign T351 = T352[5'h1f:1'h1];
  assign T352 = RouterRegFile_9_io_readData;
  assign T353 = T351[3'h4:2'h3];
  assign T354 = T351[3'h6:3'h5];
  assign T355 = T351[4'h8:3'h7];
  assign T356 = T351[4'hc:4'h9];
  assign T357 = T351[4'hd:4'hd];
  assign T358 = T351[4'he:4'he];
  assign T359 = T351[5'h1e:4'hf];
  assign T360 = T374 ? T371 : T361;
  assign T361 = T367 ? 1'h0 : T362;
  assign T362 = T363 & T301;
  assign T363 = T365 & T364;
  assign T364 = VCRouterStateManagement_9_io_currentState == 3'h4;
  assign T365 = T320 | T366;
  assign T366 = VCRouterStateManagement_9_io_currentState == 3'h4;
  assign T367 = T369 & T368;
  assign T368 = ~ RouterRegFile_9_io_readValid;
  assign T369 = T370 == 1'h1;
  assign T370 = RouterBuffer_9_io_deq_bits_x[1'h0:1'h0];
  assign T371 = T372 & T301;
  assign T372 = T365 & T373;
  assign T373 = 3'h3 <= VCRouterStateManagement_9_io_currentState;
  assign T374 = T378 & T375;
  assign T375 = T376 & RouterRegFile_9_io_readValid;
  assign T376 = T377 == 1'h1;
  assign T377 = RouterBuffer_9_io_deq_bits_x[1'h0:1'h0];
  assign T378 = T367 ^ 1'h1;
  assign T379 = io_inChannels_4_flitValid & T4;
  assign T380 = T381 & RouterRegFile_9_io_readValid;
  assign T381 = RouterRegFile_9_io_rvPipelineReg_0 ^ 1'h1;
  assign T382 = T384 & T383;
  assign T383 = VCRouterStateManagement_9_io_currentState == 3'h2;
  assign T384 = RouterRegFile_9_io_rvPipelineReg_0 & vcAllocator_io_resources_9_valid;
  assign T385 = T387 & T386;
  assign T386 = VCRouterStateManagement_9_io_currentState == 3'h3;
  assign T387 = RouterRegFile_9_io_rvPipelineReg_1 & T320;
  assign T3118 = {24'h0, T388};
  assign T388 = T389;
  assign T389 = {T393, T390};
  assign T390 = {T392, T391};
  assign T391 = {CMeshDOR_9_io_outHeadFlit_destination_0, CMeshDOR_9_io_outHeadFlit_priorityLevel};
  assign T392 = {CMeshDOR_9_io_outHeadFlit_destination_2, CMeshDOR_9_io_outHeadFlit_destination_1};
  assign T393 = {T395, T394};
  assign T394 = {CMeshDOR_9_io_outHeadFlit_vcPort, CMeshDOR_9_io_outHeadFlit_packetType};
  assign T395 = {CMeshDOR_9_io_outHeadFlit_packetID, CMeshDOR_9_io_outHeadFlit_isTail};
  assign T396 = T398 & T397;
  assign T397 = VCRouterStateManagement_9_io_currentState == 3'h4;
  assign T398 = T399 & T301;
  assign T399 = T365 & flitsAreTail_9;
  assign flitsAreTail_9 = T400;
  assign T400 = T401 & RouterBuffer_9_io_deq_valid;
  assign T401 = T402;
  assign T402 = T407 ? T405 : T403;
  assign T403 = T404[6'h25:6'h25];
  assign T404 = RouterBuffer_9_io_deq_bits_x[6'h36:1'h1];
  assign T405 = T406[4'he:4'he];
  assign T406 = RouterBuffer_9_io_deq_bits_x[5'h1f:1'h1];
  assign T407 = T408 == 1'h1;
  assign T408 = RouterBuffer_9_io_deq_bits_x[1'h0:1'h0];
  assign T409 = T410 ? T379 : 1'h0;
  assign T410 = T411 == 1'h1;
  assign T411 = io_inChannels_4_flit_x[1'h0:1'h0];
  assign T412 = T410 ? T413 : 55'h0;
  assign T413 = io_inChannels_4_flit_x;
  assign T414 = T374 ? T420 : T415;
  assign T415 = T367 ? 1'h0 : T416;
  assign T416 = T417 & RouterBuffer_9_io_deq_valid;
  assign T417 = T418 & T301;
  assign T418 = T365 & T419;
  assign T419 = VCRouterStateManagement_9_io_currentState == 3'h4;
  assign T420 = T421 & RouterBuffer_9_io_deq_valid;
  assign T421 = T422 & T301;
  assign T422 = T365 & T423;
  assign T423 = 3'h3 <= VCRouterStateManagement_9_io_currentState;
  assign T424 = T425;
  assign T425 = io_inChannels_4_flit_x;
  assign T3119 = R426[1'h0:1'h0];
  assign T3120 = reset ? 55'h0 : T427;
  assign T427 = T428 ? T3121 : R426;
  assign T3121 = {51'h0, vcAllocator_io_chosens_8};
  assign T428 = T429 & vcAllocator_io_resources_8_valid;
  assign T429 = VCRouterStateManagement_8_io_currentState == 3'h2;
  assign T430 = T431;
  assign T431 = RouterBuffer_8_io_deq_bits_x;
  assign T432 = T444 | T433;
  assign T433 = T434 == 2'h1;
  assign T434 = T443 ? VCRouterOutputStateManagement_4_io_currentState : T435;
  assign T435 = T442 ? T440 : T436;
  assign T436 = T437 ? VCRouterOutputStateManagement_1_io_currentState : VCRouterOutputStateManagement_io_currentState;
  assign T437 = T438[1'h0:1'h0];
  assign T438 = R439;
  assign T3122 = reset ? 3'h0 : CMeshDOR_8_io_result;
  assign T440 = T441 ? VCRouterOutputStateManagement_3_io_currentState : VCRouterOutputStateManagement_2_io_currentState;
  assign T441 = T438[1'h0:1'h0];
  assign T442 = T438[1'h1:1'h1];
  assign T443 = T438[2'h2:2'h2];
  assign T444 = T434 == 2'h2;
  assign T445 = T463 ? T455 : T446;
  assign T446 = T454 ? creditConsReady_4_0 : T447;
  assign T447 = T453 ? T451 : T448;
  assign T448 = T449 ? creditConsReady_1_0 : creditConsReady_0_0;
  assign T449 = T450[1'h0:1'h0];
  assign T450 = R439;
  assign T451 = T452 ? creditConsReady_3_0 : creditConsReady_2_0;
  assign T452 = T450[1'h0:1'h0];
  assign T453 = T450[1'h1:1'h1];
  assign T454 = T450[2'h2:2'h2];
  assign T455 = T462 ? creditConsReady_4_1 : T456;
  assign T456 = T461 ? T459 : T457;
  assign T457 = T458 ? creditConsReady_1_1 : creditConsReady_0_1;
  assign T458 = T450[1'h0:1'h0];
  assign T459 = T460 ? creditConsReady_3_1 : creditConsReady_2_1;
  assign T460 = T450[1'h0:1'h0];
  assign T461 = T450[1'h1:1'h1];
  assign T462 = T450[2'h2:2'h2];
  assign T463 = T3123;
  assign T3123 = R426[1'h0:1'h0];
  assign T464 = T475 & T465;
  assign T465 = T466 == 4'h8;
  assign T466 = T474 ? swAllocator_io_chosens_4 : T467;
  assign T467 = T473 ? T471 : T468;
  assign T468 = T469 ? swAllocator_io_chosens_1 : swAllocator_io_chosens_0;
  assign T469 = T470[1'h0:1'h0];
  assign T470 = R439;
  assign T471 = T472 ? swAllocator_io_chosens_3 : swAllocator_io_chosens_2;
  assign T472 = T470[1'h0:1'h0];
  assign T473 = T470[1'h1:1'h1];
  assign T474 = T470[2'h2:2'h2];
  assign T475 = T483 ? swAllocator_io_requests_4_8_grant : T476;
  assign T476 = T482 ? T480 : T477;
  assign T477 = T478 ? swAllocator_io_requests_1_8_grant : swAllocator_io_requests_0_8_grant;
  assign T478 = T479[1'h0:1'h0];
  assign T479 = R439;
  assign T480 = T481 ? swAllocator_io_requests_3_8_grant : swAllocator_io_requests_2_8_grant;
  assign T481 = T479[1'h0:1'h0];
  assign T482 = T479[1'h1:1'h1];
  assign T483 = T479[2'h2:2'h2];
  assign T484 = RouterBuffer_8_io_deq_valid & T485;
  assign T485 = T486;
  assign T486 = T491 ? T489 : T487;
  assign T487 = T488[6'h25:6'h25];
  assign T488 = RouterBuffer_8_io_deq_bits_x[6'h36:1'h1];
  assign T489 = T490[4'he:4'he];
  assign T490 = RouterBuffer_8_io_deq_bits_x[5'h1f:1'h1];
  assign T491 = T492 == 1'h1;
  assign T492 = RouterBuffer_8_io_deq_bits_x[1'h0:1'h0];
  assign T3124 = reset ? 1'h0 : RouterBuffer_8_io_deq_valid;
  assign T494 = T495[2'h2:1'h0];
  assign T495 = T496[5'h1f:1'h1];
  assign T496 = RouterRegFile_8_io_readData;
  assign T497 = T495[3'h4:2'h3];
  assign T498 = T495[3'h6:3'h5];
  assign T499 = T495[4'h8:3'h7];
  assign T500 = T495[4'hc:4'h9];
  assign T501 = T495[4'hd:4'hd];
  assign T502 = T495[4'he:4'he];
  assign T503 = T495[5'h1e:4'hf];
  assign T504 = T518 ? T515 : T505;
  assign T505 = T511 ? 1'h0 : T506;
  assign T506 = T507 & T445;
  assign T507 = T509 & T508;
  assign T508 = VCRouterStateManagement_8_io_currentState == 3'h4;
  assign T509 = T464 | T510;
  assign T510 = VCRouterStateManagement_8_io_currentState == 3'h4;
  assign T511 = T513 & T512;
  assign T512 = ~ RouterRegFile_8_io_readValid;
  assign T513 = T514 == 1'h1;
  assign T514 = RouterBuffer_8_io_deq_bits_x[1'h0:1'h0];
  assign T515 = T516 & T445;
  assign T516 = T509 & T517;
  assign T517 = 3'h3 <= VCRouterStateManagement_8_io_currentState;
  assign T518 = T522 & T519;
  assign T519 = T520 & RouterRegFile_8_io_readValid;
  assign T520 = T521 == 1'h1;
  assign T521 = RouterBuffer_8_io_deq_bits_x[1'h0:1'h0];
  assign T522 = T511 ^ 1'h1;
  assign T523 = io_inChannels_4_flitValid & T26;
  assign T524 = T525 & RouterRegFile_8_io_readValid;
  assign T525 = RouterRegFile_8_io_rvPipelineReg_0 ^ 1'h1;
  assign T526 = T528 & T527;
  assign T527 = VCRouterStateManagement_8_io_currentState == 3'h2;
  assign T528 = RouterRegFile_8_io_rvPipelineReg_0 & vcAllocator_io_resources_8_valid;
  assign T529 = T531 & T530;
  assign T530 = VCRouterStateManagement_8_io_currentState == 3'h3;
  assign T531 = RouterRegFile_8_io_rvPipelineReg_1 & T464;
  assign T3125 = {24'h0, T532};
  assign T532 = T533;
  assign T533 = {T537, T534};
  assign T534 = {T536, T535};
  assign T535 = {CMeshDOR_8_io_outHeadFlit_destination_0, CMeshDOR_8_io_outHeadFlit_priorityLevel};
  assign T536 = {CMeshDOR_8_io_outHeadFlit_destination_2, CMeshDOR_8_io_outHeadFlit_destination_1};
  assign T537 = {T539, T538};
  assign T538 = {CMeshDOR_8_io_outHeadFlit_vcPort, CMeshDOR_8_io_outHeadFlit_packetType};
  assign T539 = {CMeshDOR_8_io_outHeadFlit_packetID, CMeshDOR_8_io_outHeadFlit_isTail};
  assign T540 = T542 & T541;
  assign T541 = VCRouterStateManagement_8_io_currentState == 3'h4;
  assign T542 = T543 & T445;
  assign T543 = T509 & flitsAreTail_8;
  assign flitsAreTail_8 = T544;
  assign T544 = T545 & RouterBuffer_8_io_deq_valid;
  assign T545 = T546;
  assign T546 = T551 ? T549 : T547;
  assign T547 = T548[6'h25:6'h25];
  assign T548 = RouterBuffer_8_io_deq_bits_x[6'h36:1'h1];
  assign T549 = T550[4'he:4'he];
  assign T550 = RouterBuffer_8_io_deq_bits_x[5'h1f:1'h1];
  assign T551 = T552 == 1'h1;
  assign T552 = RouterBuffer_8_io_deq_bits_x[1'h0:1'h0];
  assign T553 = T554 ? T523 : 1'h0;
  assign T554 = T555 == 1'h1;
  assign T555 = io_inChannels_4_flit_x[1'h0:1'h0];
  assign T556 = T554 ? T557 : 55'h0;
  assign T557 = io_inChannels_4_flit_x;
  assign T558 = T518 ? T564 : T559;
  assign T559 = T511 ? 1'h0 : T560;
  assign T560 = T561 & RouterBuffer_8_io_deq_valid;
  assign T561 = T562 & T445;
  assign T562 = T509 & T563;
  assign T563 = VCRouterStateManagement_8_io_currentState == 3'h4;
  assign T564 = T565 & RouterBuffer_8_io_deq_valid;
  assign T565 = T566 & T445;
  assign T566 = T509 & T567;
  assign T567 = 3'h3 <= VCRouterStateManagement_8_io_currentState;
  assign T568 = T569;
  assign T569 = io_inChannels_3_flit_x;
  assign T3126 = R570[1'h0:1'h0];
  assign T3127 = reset ? 55'h0 : T571;
  assign T571 = T572 ? T3128 : R570;
  assign T3128 = {51'h0, vcAllocator_io_chosens_7};
  assign T572 = T573 & vcAllocator_io_resources_7_valid;
  assign T573 = VCRouterStateManagement_7_io_currentState == 3'h2;
  assign T574 = T575;
  assign T575 = RouterBuffer_7_io_deq_bits_x;
  assign T576 = T588 | T577;
  assign T577 = T578 == 2'h1;
  assign T578 = T587 ? VCRouterOutputStateManagement_4_io_currentState : T579;
  assign T579 = T586 ? T584 : T580;
  assign T580 = T581 ? VCRouterOutputStateManagement_1_io_currentState : VCRouterOutputStateManagement_io_currentState;
  assign T581 = T582[1'h0:1'h0];
  assign T582 = R583;
  assign T3129 = reset ? 3'h0 : CMeshDOR_7_io_result;
  assign T584 = T585 ? VCRouterOutputStateManagement_3_io_currentState : VCRouterOutputStateManagement_2_io_currentState;
  assign T585 = T582[1'h0:1'h0];
  assign T586 = T582[1'h1:1'h1];
  assign T587 = T582[2'h2:2'h2];
  assign T588 = T578 == 2'h2;
  assign T589 = T607 ? T599 : T590;
  assign T590 = T598 ? creditConsReady_4_0 : T591;
  assign T591 = T597 ? T595 : T592;
  assign T592 = T593 ? creditConsReady_1_0 : creditConsReady_0_0;
  assign T593 = T594[1'h0:1'h0];
  assign T594 = R583;
  assign T595 = T596 ? creditConsReady_3_0 : creditConsReady_2_0;
  assign T596 = T594[1'h0:1'h0];
  assign T597 = T594[1'h1:1'h1];
  assign T598 = T594[2'h2:2'h2];
  assign T599 = T606 ? creditConsReady_4_1 : T600;
  assign T600 = T605 ? T603 : T601;
  assign T601 = T602 ? creditConsReady_1_1 : creditConsReady_0_1;
  assign T602 = T594[1'h0:1'h0];
  assign T603 = T604 ? creditConsReady_3_1 : creditConsReady_2_1;
  assign T604 = T594[1'h0:1'h0];
  assign T605 = T594[1'h1:1'h1];
  assign T606 = T594[2'h2:2'h2];
  assign T607 = T3130;
  assign T3130 = R570[1'h0:1'h0];
  assign T608 = T619 & T609;
  assign T609 = T610 == 4'h7;
  assign T610 = T618 ? swAllocator_io_chosens_4 : T611;
  assign T611 = T617 ? T615 : T612;
  assign T612 = T613 ? swAllocator_io_chosens_1 : swAllocator_io_chosens_0;
  assign T613 = T614[1'h0:1'h0];
  assign T614 = R583;
  assign T615 = T616 ? swAllocator_io_chosens_3 : swAllocator_io_chosens_2;
  assign T616 = T614[1'h0:1'h0];
  assign T617 = T614[1'h1:1'h1];
  assign T618 = T614[2'h2:2'h2];
  assign T619 = T627 ? swAllocator_io_requests_4_7_grant : T620;
  assign T620 = T626 ? T624 : T621;
  assign T621 = T622 ? swAllocator_io_requests_1_7_grant : swAllocator_io_requests_0_7_grant;
  assign T622 = T623[1'h0:1'h0];
  assign T623 = R583;
  assign T624 = T625 ? swAllocator_io_requests_3_7_grant : swAllocator_io_requests_2_7_grant;
  assign T625 = T623[1'h0:1'h0];
  assign T626 = T623[1'h1:1'h1];
  assign T627 = T623[2'h2:2'h2];
  assign T628 = RouterBuffer_7_io_deq_valid & T629;
  assign T629 = T630;
  assign T630 = T635 ? T633 : T631;
  assign T631 = T632[6'h25:6'h25];
  assign T632 = RouterBuffer_7_io_deq_bits_x[6'h36:1'h1];
  assign T633 = T634[4'he:4'he];
  assign T634 = RouterBuffer_7_io_deq_bits_x[5'h1f:1'h1];
  assign T635 = T636 == 1'h1;
  assign T636 = RouterBuffer_7_io_deq_bits_x[1'h0:1'h0];
  assign T3131 = reset ? 1'h0 : RouterBuffer_7_io_deq_valid;
  assign T638 = T639[2'h2:1'h0];
  assign T639 = T640[5'h1f:1'h1];
  assign T640 = RouterRegFile_7_io_readData;
  assign T641 = T639[3'h4:2'h3];
  assign T642 = T639[3'h6:3'h5];
  assign T643 = T639[4'h8:3'h7];
  assign T644 = T639[4'hc:4'h9];
  assign T645 = T639[4'hd:4'hd];
  assign T646 = T639[4'he:4'he];
  assign T647 = T639[5'h1e:4'hf];
  assign T648 = T662 ? T659 : T649;
  assign T649 = T655 ? 1'h0 : T650;
  assign T650 = T651 & T589;
  assign T651 = T653 & T652;
  assign T652 = VCRouterStateManagement_7_io_currentState == 3'h4;
  assign T653 = T608 | T654;
  assign T654 = VCRouterStateManagement_7_io_currentState == 3'h4;
  assign T655 = T657 & T656;
  assign T656 = ~ RouterRegFile_7_io_readValid;
  assign T657 = T658 == 1'h1;
  assign T658 = RouterBuffer_7_io_deq_bits_x[1'h0:1'h0];
  assign T659 = T660 & T589;
  assign T660 = T653 & T661;
  assign T661 = 3'h3 <= VCRouterStateManagement_7_io_currentState;
  assign T662 = T666 & T663;
  assign T663 = T664 & RouterRegFile_7_io_readValid;
  assign T664 = T665 == 1'h1;
  assign T665 = RouterBuffer_7_io_deq_bits_x[1'h0:1'h0];
  assign T666 = T655 ^ 1'h1;
  assign T667 = io_inChannels_3_flitValid & T48;
  assign T668 = T669 & RouterRegFile_7_io_readValid;
  assign T669 = RouterRegFile_7_io_rvPipelineReg_0 ^ 1'h1;
  assign T670 = T672 & T671;
  assign T671 = VCRouterStateManagement_7_io_currentState == 3'h2;
  assign T672 = RouterRegFile_7_io_rvPipelineReg_0 & vcAllocator_io_resources_7_valid;
  assign T673 = T675 & T674;
  assign T674 = VCRouterStateManagement_7_io_currentState == 3'h3;
  assign T675 = RouterRegFile_7_io_rvPipelineReg_1 & T608;
  assign T3132 = {24'h0, T676};
  assign T676 = T677;
  assign T677 = {T681, T678};
  assign T678 = {T680, T679};
  assign T679 = {CMeshDOR_7_io_outHeadFlit_destination_0, CMeshDOR_7_io_outHeadFlit_priorityLevel};
  assign T680 = {CMeshDOR_7_io_outHeadFlit_destination_2, CMeshDOR_7_io_outHeadFlit_destination_1};
  assign T681 = {T683, T682};
  assign T682 = {CMeshDOR_7_io_outHeadFlit_vcPort, CMeshDOR_7_io_outHeadFlit_packetType};
  assign T683 = {CMeshDOR_7_io_outHeadFlit_packetID, CMeshDOR_7_io_outHeadFlit_isTail};
  assign T684 = T686 & T685;
  assign T685 = VCRouterStateManagement_7_io_currentState == 3'h4;
  assign T686 = T687 & T589;
  assign T687 = T653 & flitsAreTail_7;
  assign flitsAreTail_7 = T688;
  assign T688 = T689 & RouterBuffer_7_io_deq_valid;
  assign T689 = T690;
  assign T690 = T695 ? T693 : T691;
  assign T691 = T692[6'h25:6'h25];
  assign T692 = RouterBuffer_7_io_deq_bits_x[6'h36:1'h1];
  assign T693 = T694[4'he:4'he];
  assign T694 = RouterBuffer_7_io_deq_bits_x[5'h1f:1'h1];
  assign T695 = T696 == 1'h1;
  assign T696 = RouterBuffer_7_io_deq_bits_x[1'h0:1'h0];
  assign T697 = T698 ? T667 : 1'h0;
  assign T698 = T699 == 1'h1;
  assign T699 = io_inChannels_3_flit_x[1'h0:1'h0];
  assign T700 = T698 ? T701 : 55'h0;
  assign T701 = io_inChannels_3_flit_x;
  assign T702 = T662 ? T708 : T703;
  assign T703 = T655 ? 1'h0 : T704;
  assign T704 = T705 & RouterBuffer_7_io_deq_valid;
  assign T705 = T706 & T589;
  assign T706 = T653 & T707;
  assign T707 = VCRouterStateManagement_7_io_currentState == 3'h4;
  assign T708 = T709 & RouterBuffer_7_io_deq_valid;
  assign T709 = T710 & T589;
  assign T710 = T653 & T711;
  assign T711 = 3'h3 <= VCRouterStateManagement_7_io_currentState;
  assign T712 = T713;
  assign T713 = io_inChannels_3_flit_x;
  assign T3133 = R714[1'h0:1'h0];
  assign T3134 = reset ? 55'h0 : T715;
  assign T715 = T716 ? T3135 : R714;
  assign T3135 = {51'h0, vcAllocator_io_chosens_6};
  assign T716 = T717 & vcAllocator_io_resources_6_valid;
  assign T717 = VCRouterStateManagement_6_io_currentState == 3'h2;
  assign T718 = T719;
  assign T719 = RouterBuffer_6_io_deq_bits_x;
  assign T720 = T732 | T721;
  assign T721 = T722 == 2'h1;
  assign T722 = T731 ? VCRouterOutputStateManagement_4_io_currentState : T723;
  assign T723 = T730 ? T728 : T724;
  assign T724 = T725 ? VCRouterOutputStateManagement_1_io_currentState : VCRouterOutputStateManagement_io_currentState;
  assign T725 = T726[1'h0:1'h0];
  assign T726 = R727;
  assign T3136 = reset ? 3'h0 : CMeshDOR_6_io_result;
  assign T728 = T729 ? VCRouterOutputStateManagement_3_io_currentState : VCRouterOutputStateManagement_2_io_currentState;
  assign T729 = T726[1'h0:1'h0];
  assign T730 = T726[1'h1:1'h1];
  assign T731 = T726[2'h2:2'h2];
  assign T732 = T722 == 2'h2;
  assign T733 = T751 ? T743 : T734;
  assign T734 = T742 ? creditConsReady_4_0 : T735;
  assign T735 = T741 ? T739 : T736;
  assign T736 = T737 ? creditConsReady_1_0 : creditConsReady_0_0;
  assign T737 = T738[1'h0:1'h0];
  assign T738 = R727;
  assign T739 = T740 ? creditConsReady_3_0 : creditConsReady_2_0;
  assign T740 = T738[1'h0:1'h0];
  assign T741 = T738[1'h1:1'h1];
  assign T742 = T738[2'h2:2'h2];
  assign T743 = T750 ? creditConsReady_4_1 : T744;
  assign T744 = T749 ? T747 : T745;
  assign T745 = T746 ? creditConsReady_1_1 : creditConsReady_0_1;
  assign T746 = T738[1'h0:1'h0];
  assign T747 = T748 ? creditConsReady_3_1 : creditConsReady_2_1;
  assign T748 = T738[1'h0:1'h0];
  assign T749 = T738[1'h1:1'h1];
  assign T750 = T738[2'h2:2'h2];
  assign T751 = T3137;
  assign T3137 = R714[1'h0:1'h0];
  assign T752 = T763 & T753;
  assign T753 = T754 == 4'h6;
  assign T754 = T762 ? swAllocator_io_chosens_4 : T755;
  assign T755 = T761 ? T759 : T756;
  assign T756 = T757 ? swAllocator_io_chosens_1 : swAllocator_io_chosens_0;
  assign T757 = T758[1'h0:1'h0];
  assign T758 = R727;
  assign T759 = T760 ? swAllocator_io_chosens_3 : swAllocator_io_chosens_2;
  assign T760 = T758[1'h0:1'h0];
  assign T761 = T758[1'h1:1'h1];
  assign T762 = T758[2'h2:2'h2];
  assign T763 = T771 ? swAllocator_io_requests_4_6_grant : T764;
  assign T764 = T770 ? T768 : T765;
  assign T765 = T766 ? swAllocator_io_requests_1_6_grant : swAllocator_io_requests_0_6_grant;
  assign T766 = T767[1'h0:1'h0];
  assign T767 = R727;
  assign T768 = T769 ? swAllocator_io_requests_3_6_grant : swAllocator_io_requests_2_6_grant;
  assign T769 = T767[1'h0:1'h0];
  assign T770 = T767[1'h1:1'h1];
  assign T771 = T767[2'h2:2'h2];
  assign T772 = RouterBuffer_6_io_deq_valid & T773;
  assign T773 = T774;
  assign T774 = T779 ? T777 : T775;
  assign T775 = T776[6'h25:6'h25];
  assign T776 = RouterBuffer_6_io_deq_bits_x[6'h36:1'h1];
  assign T777 = T778[4'he:4'he];
  assign T778 = RouterBuffer_6_io_deq_bits_x[5'h1f:1'h1];
  assign T779 = T780 == 1'h1;
  assign T780 = RouterBuffer_6_io_deq_bits_x[1'h0:1'h0];
  assign T3138 = reset ? 1'h0 : RouterBuffer_6_io_deq_valid;
  assign T782 = T783[2'h2:1'h0];
  assign T783 = T784[5'h1f:1'h1];
  assign T784 = RouterRegFile_6_io_readData;
  assign T785 = T783[3'h4:2'h3];
  assign T786 = T783[3'h6:3'h5];
  assign T787 = T783[4'h8:3'h7];
  assign T788 = T783[4'hc:4'h9];
  assign T789 = T783[4'hd:4'hd];
  assign T790 = T783[4'he:4'he];
  assign T791 = T783[5'h1e:4'hf];
  assign T792 = T806 ? T803 : T793;
  assign T793 = T799 ? 1'h0 : T794;
  assign T794 = T795 & T733;
  assign T795 = T797 & T796;
  assign T796 = VCRouterStateManagement_6_io_currentState == 3'h4;
  assign T797 = T752 | T798;
  assign T798 = VCRouterStateManagement_6_io_currentState == 3'h4;
  assign T799 = T801 & T800;
  assign T800 = ~ RouterRegFile_6_io_readValid;
  assign T801 = T802 == 1'h1;
  assign T802 = RouterBuffer_6_io_deq_bits_x[1'h0:1'h0];
  assign T803 = T804 & T733;
  assign T804 = T797 & T805;
  assign T805 = 3'h3 <= VCRouterStateManagement_6_io_currentState;
  assign T806 = T810 & T807;
  assign T807 = T808 & RouterRegFile_6_io_readValid;
  assign T808 = T809 == 1'h1;
  assign T809 = RouterBuffer_6_io_deq_bits_x[1'h0:1'h0];
  assign T810 = T799 ^ 1'h1;
  assign T811 = io_inChannels_3_flitValid & T70;
  assign T812 = T813 & RouterRegFile_6_io_readValid;
  assign T813 = RouterRegFile_6_io_rvPipelineReg_0 ^ 1'h1;
  assign T814 = T816 & T815;
  assign T815 = VCRouterStateManagement_6_io_currentState == 3'h2;
  assign T816 = RouterRegFile_6_io_rvPipelineReg_0 & vcAllocator_io_resources_6_valid;
  assign T817 = T819 & T818;
  assign T818 = VCRouterStateManagement_6_io_currentState == 3'h3;
  assign T819 = RouterRegFile_6_io_rvPipelineReg_1 & T752;
  assign T3139 = {24'h0, T820};
  assign T820 = T821;
  assign T821 = {T825, T822};
  assign T822 = {T824, T823};
  assign T823 = {CMeshDOR_6_io_outHeadFlit_destination_0, CMeshDOR_6_io_outHeadFlit_priorityLevel};
  assign T824 = {CMeshDOR_6_io_outHeadFlit_destination_2, CMeshDOR_6_io_outHeadFlit_destination_1};
  assign T825 = {T827, T826};
  assign T826 = {CMeshDOR_6_io_outHeadFlit_vcPort, CMeshDOR_6_io_outHeadFlit_packetType};
  assign T827 = {CMeshDOR_6_io_outHeadFlit_packetID, CMeshDOR_6_io_outHeadFlit_isTail};
  assign T828 = T830 & T829;
  assign T829 = VCRouterStateManagement_6_io_currentState == 3'h4;
  assign T830 = T831 & T733;
  assign T831 = T797 & flitsAreTail_6;
  assign flitsAreTail_6 = T832;
  assign T832 = T833 & RouterBuffer_6_io_deq_valid;
  assign T833 = T834;
  assign T834 = T839 ? T837 : T835;
  assign T835 = T836[6'h25:6'h25];
  assign T836 = RouterBuffer_6_io_deq_bits_x[6'h36:1'h1];
  assign T837 = T838[4'he:4'he];
  assign T838 = RouterBuffer_6_io_deq_bits_x[5'h1f:1'h1];
  assign T839 = T840 == 1'h1;
  assign T840 = RouterBuffer_6_io_deq_bits_x[1'h0:1'h0];
  assign T841 = T842 ? T811 : 1'h0;
  assign T842 = T843 == 1'h1;
  assign T843 = io_inChannels_3_flit_x[1'h0:1'h0];
  assign T844 = T842 ? T845 : 55'h0;
  assign T845 = io_inChannels_3_flit_x;
  assign T846 = T806 ? T852 : T847;
  assign T847 = T799 ? 1'h0 : T848;
  assign T848 = T849 & RouterBuffer_6_io_deq_valid;
  assign T849 = T850 & T733;
  assign T850 = T797 & T851;
  assign T851 = VCRouterStateManagement_6_io_currentState == 3'h4;
  assign T852 = T853 & RouterBuffer_6_io_deq_valid;
  assign T853 = T854 & T733;
  assign T854 = T797 & T855;
  assign T855 = 3'h3 <= VCRouterStateManagement_6_io_currentState;
  assign T856 = T857;
  assign T857 = io_inChannels_2_flit_x;
  assign T3140 = R858[1'h0:1'h0];
  assign T3141 = reset ? 55'h0 : T859;
  assign T859 = T860 ? T3142 : R858;
  assign T3142 = {51'h0, vcAllocator_io_chosens_5};
  assign T860 = T861 & vcAllocator_io_resources_5_valid;
  assign T861 = VCRouterStateManagement_5_io_currentState == 3'h2;
  assign T862 = T863;
  assign T863 = RouterBuffer_5_io_deq_bits_x;
  assign T864 = T876 | T865;
  assign T865 = T866 == 2'h1;
  assign T866 = T875 ? VCRouterOutputStateManagement_4_io_currentState : T867;
  assign T867 = T874 ? T872 : T868;
  assign T868 = T869 ? VCRouterOutputStateManagement_1_io_currentState : VCRouterOutputStateManagement_io_currentState;
  assign T869 = T870[1'h0:1'h0];
  assign T870 = R871;
  assign T3143 = reset ? 3'h0 : CMeshDOR_5_io_result;
  assign T872 = T873 ? VCRouterOutputStateManagement_3_io_currentState : VCRouterOutputStateManagement_2_io_currentState;
  assign T873 = T870[1'h0:1'h0];
  assign T874 = T870[1'h1:1'h1];
  assign T875 = T870[2'h2:2'h2];
  assign T876 = T866 == 2'h2;
  assign T877 = T895 ? T887 : T878;
  assign T878 = T886 ? creditConsReady_4_0 : T879;
  assign T879 = T885 ? T883 : T880;
  assign T880 = T881 ? creditConsReady_1_0 : creditConsReady_0_0;
  assign T881 = T882[1'h0:1'h0];
  assign T882 = R871;
  assign T883 = T884 ? creditConsReady_3_0 : creditConsReady_2_0;
  assign T884 = T882[1'h0:1'h0];
  assign T885 = T882[1'h1:1'h1];
  assign T886 = T882[2'h2:2'h2];
  assign T887 = T894 ? creditConsReady_4_1 : T888;
  assign T888 = T893 ? T891 : T889;
  assign T889 = T890 ? creditConsReady_1_1 : creditConsReady_0_1;
  assign T890 = T882[1'h0:1'h0];
  assign T891 = T892 ? creditConsReady_3_1 : creditConsReady_2_1;
  assign T892 = T882[1'h0:1'h0];
  assign T893 = T882[1'h1:1'h1];
  assign T894 = T882[2'h2:2'h2];
  assign T895 = T3144;
  assign T3144 = R858[1'h0:1'h0];
  assign T896 = T907 & T897;
  assign T897 = T898 == 4'h5;
  assign T898 = T906 ? swAllocator_io_chosens_4 : T899;
  assign T899 = T905 ? T903 : T900;
  assign T900 = T901 ? swAllocator_io_chosens_1 : swAllocator_io_chosens_0;
  assign T901 = T902[1'h0:1'h0];
  assign T902 = R871;
  assign T903 = T904 ? swAllocator_io_chosens_3 : swAllocator_io_chosens_2;
  assign T904 = T902[1'h0:1'h0];
  assign T905 = T902[1'h1:1'h1];
  assign T906 = T902[2'h2:2'h2];
  assign T907 = T915 ? swAllocator_io_requests_4_5_grant : T908;
  assign T908 = T914 ? T912 : T909;
  assign T909 = T910 ? swAllocator_io_requests_1_5_grant : swAllocator_io_requests_0_5_grant;
  assign T910 = T911[1'h0:1'h0];
  assign T911 = R871;
  assign T912 = T913 ? swAllocator_io_requests_3_5_grant : swAllocator_io_requests_2_5_grant;
  assign T913 = T911[1'h0:1'h0];
  assign T914 = T911[1'h1:1'h1];
  assign T915 = T911[2'h2:2'h2];
  assign T916 = RouterBuffer_5_io_deq_valid & T917;
  assign T917 = T918;
  assign T918 = T923 ? T921 : T919;
  assign T919 = T920[6'h25:6'h25];
  assign T920 = RouterBuffer_5_io_deq_bits_x[6'h36:1'h1];
  assign T921 = T922[4'he:4'he];
  assign T922 = RouterBuffer_5_io_deq_bits_x[5'h1f:1'h1];
  assign T923 = T924 == 1'h1;
  assign T924 = RouterBuffer_5_io_deq_bits_x[1'h0:1'h0];
  assign T3145 = reset ? 1'h0 : RouterBuffer_5_io_deq_valid;
  assign T926 = T927[2'h2:1'h0];
  assign T927 = T928[5'h1f:1'h1];
  assign T928 = RouterRegFile_5_io_readData;
  assign T929 = T927[3'h4:2'h3];
  assign T930 = T927[3'h6:3'h5];
  assign T931 = T927[4'h8:3'h7];
  assign T932 = T927[4'hc:4'h9];
  assign T933 = T927[4'hd:4'hd];
  assign T934 = T927[4'he:4'he];
  assign T935 = T927[5'h1e:4'hf];
  assign T936 = T950 ? T947 : T937;
  assign T937 = T943 ? 1'h0 : T938;
  assign T938 = T939 & T877;
  assign T939 = T941 & T940;
  assign T940 = VCRouterStateManagement_5_io_currentState == 3'h4;
  assign T941 = T896 | T942;
  assign T942 = VCRouterStateManagement_5_io_currentState == 3'h4;
  assign T943 = T945 & T944;
  assign T944 = ~ RouterRegFile_5_io_readValid;
  assign T945 = T946 == 1'h1;
  assign T946 = RouterBuffer_5_io_deq_bits_x[1'h0:1'h0];
  assign T947 = T948 & T877;
  assign T948 = T941 & T949;
  assign T949 = 3'h3 <= VCRouterStateManagement_5_io_currentState;
  assign T950 = T954 & T951;
  assign T951 = T952 & RouterRegFile_5_io_readValid;
  assign T952 = T953 == 1'h1;
  assign T953 = RouterBuffer_5_io_deq_bits_x[1'h0:1'h0];
  assign T954 = T943 ^ 1'h1;
  assign T955 = io_inChannels_2_flitValid & T92;
  assign T956 = T957 & RouterRegFile_5_io_readValid;
  assign T957 = RouterRegFile_5_io_rvPipelineReg_0 ^ 1'h1;
  assign T958 = T960 & T959;
  assign T959 = VCRouterStateManagement_5_io_currentState == 3'h2;
  assign T960 = RouterRegFile_5_io_rvPipelineReg_0 & vcAllocator_io_resources_5_valid;
  assign T961 = T963 & T962;
  assign T962 = VCRouterStateManagement_5_io_currentState == 3'h3;
  assign T963 = RouterRegFile_5_io_rvPipelineReg_1 & T896;
  assign T3146 = {24'h0, T964};
  assign T964 = T965;
  assign T965 = {T969, T966};
  assign T966 = {T968, T967};
  assign T967 = {CMeshDOR_5_io_outHeadFlit_destination_0, CMeshDOR_5_io_outHeadFlit_priorityLevel};
  assign T968 = {CMeshDOR_5_io_outHeadFlit_destination_2, CMeshDOR_5_io_outHeadFlit_destination_1};
  assign T969 = {T971, T970};
  assign T970 = {CMeshDOR_5_io_outHeadFlit_vcPort, CMeshDOR_5_io_outHeadFlit_packetType};
  assign T971 = {CMeshDOR_5_io_outHeadFlit_packetID, CMeshDOR_5_io_outHeadFlit_isTail};
  assign T972 = T974 & T973;
  assign T973 = VCRouterStateManagement_5_io_currentState == 3'h4;
  assign T974 = T975 & T877;
  assign T975 = T941 & flitsAreTail_5;
  assign flitsAreTail_5 = T976;
  assign T976 = T977 & RouterBuffer_5_io_deq_valid;
  assign T977 = T978;
  assign T978 = T983 ? T981 : T979;
  assign T979 = T980[6'h25:6'h25];
  assign T980 = RouterBuffer_5_io_deq_bits_x[6'h36:1'h1];
  assign T981 = T982[4'he:4'he];
  assign T982 = RouterBuffer_5_io_deq_bits_x[5'h1f:1'h1];
  assign T983 = T984 == 1'h1;
  assign T984 = RouterBuffer_5_io_deq_bits_x[1'h0:1'h0];
  assign T985 = T986 ? T955 : 1'h0;
  assign T986 = T987 == 1'h1;
  assign T987 = io_inChannels_2_flit_x[1'h0:1'h0];
  assign T988 = T986 ? T989 : 55'h0;
  assign T989 = io_inChannels_2_flit_x;
  assign T990 = T950 ? T996 : T991;
  assign T991 = T943 ? 1'h0 : T992;
  assign T992 = T993 & RouterBuffer_5_io_deq_valid;
  assign T993 = T994 & T877;
  assign T994 = T941 & T995;
  assign T995 = VCRouterStateManagement_5_io_currentState == 3'h4;
  assign T996 = T997 & RouterBuffer_5_io_deq_valid;
  assign T997 = T998 & T877;
  assign T998 = T941 & T999;
  assign T999 = 3'h3 <= VCRouterStateManagement_5_io_currentState;
  assign T1000 = T1001;
  assign T1001 = io_inChannels_2_flit_x;
  assign T3147 = R1002[1'h0:1'h0];
  assign T3148 = reset ? 55'h0 : T1003;
  assign T1003 = T1004 ? T3149 : R1002;
  assign T3149 = {51'h0, vcAllocator_io_chosens_4};
  assign T1004 = T1005 & vcAllocator_io_resources_4_valid;
  assign T1005 = VCRouterStateManagement_4_io_currentState == 3'h2;
  assign T1006 = T1007;
  assign T1007 = RouterBuffer_4_io_deq_bits_x;
  assign T1008 = T1020 | T1009;
  assign T1009 = T1010 == 2'h1;
  assign T1010 = T1019 ? VCRouterOutputStateManagement_4_io_currentState : T1011;
  assign T1011 = T1018 ? T1016 : T1012;
  assign T1012 = T1013 ? VCRouterOutputStateManagement_1_io_currentState : VCRouterOutputStateManagement_io_currentState;
  assign T1013 = T1014[1'h0:1'h0];
  assign T1014 = R1015;
  assign T3150 = reset ? 3'h0 : CMeshDOR_4_io_result;
  assign T1016 = T1017 ? VCRouterOutputStateManagement_3_io_currentState : VCRouterOutputStateManagement_2_io_currentState;
  assign T1017 = T1014[1'h0:1'h0];
  assign T1018 = T1014[1'h1:1'h1];
  assign T1019 = T1014[2'h2:2'h2];
  assign T1020 = T1010 == 2'h2;
  assign T1021 = T1039 ? T1031 : T1022;
  assign T1022 = T1030 ? creditConsReady_4_0 : T1023;
  assign T1023 = T1029 ? T1027 : T1024;
  assign T1024 = T1025 ? creditConsReady_1_0 : creditConsReady_0_0;
  assign T1025 = T1026[1'h0:1'h0];
  assign T1026 = R1015;
  assign T1027 = T1028 ? creditConsReady_3_0 : creditConsReady_2_0;
  assign T1028 = T1026[1'h0:1'h0];
  assign T1029 = T1026[1'h1:1'h1];
  assign T1030 = T1026[2'h2:2'h2];
  assign T1031 = T1038 ? creditConsReady_4_1 : T1032;
  assign T1032 = T1037 ? T1035 : T1033;
  assign T1033 = T1034 ? creditConsReady_1_1 : creditConsReady_0_1;
  assign T1034 = T1026[1'h0:1'h0];
  assign T1035 = T1036 ? creditConsReady_3_1 : creditConsReady_2_1;
  assign T1036 = T1026[1'h0:1'h0];
  assign T1037 = T1026[1'h1:1'h1];
  assign T1038 = T1026[2'h2:2'h2];
  assign T1039 = T3151;
  assign T3151 = R1002[1'h0:1'h0];
  assign T1040 = T1051 & T1041;
  assign T1041 = T1042 == 4'h4;
  assign T1042 = T1050 ? swAllocator_io_chosens_4 : T1043;
  assign T1043 = T1049 ? T1047 : T1044;
  assign T1044 = T1045 ? swAllocator_io_chosens_1 : swAllocator_io_chosens_0;
  assign T1045 = T1046[1'h0:1'h0];
  assign T1046 = R1015;
  assign T1047 = T1048 ? swAllocator_io_chosens_3 : swAllocator_io_chosens_2;
  assign T1048 = T1046[1'h0:1'h0];
  assign T1049 = T1046[1'h1:1'h1];
  assign T1050 = T1046[2'h2:2'h2];
  assign T1051 = T1059 ? swAllocator_io_requests_4_4_grant : T1052;
  assign T1052 = T1058 ? T1056 : T1053;
  assign T1053 = T1054 ? swAllocator_io_requests_1_4_grant : swAllocator_io_requests_0_4_grant;
  assign T1054 = T1055[1'h0:1'h0];
  assign T1055 = R1015;
  assign T1056 = T1057 ? swAllocator_io_requests_3_4_grant : swAllocator_io_requests_2_4_grant;
  assign T1057 = T1055[1'h0:1'h0];
  assign T1058 = T1055[1'h1:1'h1];
  assign T1059 = T1055[2'h2:2'h2];
  assign T1060 = RouterBuffer_4_io_deq_valid & T1061;
  assign T1061 = T1062;
  assign T1062 = T1067 ? T1065 : T1063;
  assign T1063 = T1064[6'h25:6'h25];
  assign T1064 = RouterBuffer_4_io_deq_bits_x[6'h36:1'h1];
  assign T1065 = T1066[4'he:4'he];
  assign T1066 = RouterBuffer_4_io_deq_bits_x[5'h1f:1'h1];
  assign T1067 = T1068 == 1'h1;
  assign T1068 = RouterBuffer_4_io_deq_bits_x[1'h0:1'h0];
  assign T3152 = reset ? 1'h0 : RouterBuffer_4_io_deq_valid;
  assign T1070 = T1071[2'h2:1'h0];
  assign T1071 = T1072[5'h1f:1'h1];
  assign T1072 = RouterRegFile_4_io_readData;
  assign T1073 = T1071[3'h4:2'h3];
  assign T1074 = T1071[3'h6:3'h5];
  assign T1075 = T1071[4'h8:3'h7];
  assign T1076 = T1071[4'hc:4'h9];
  assign T1077 = T1071[4'hd:4'hd];
  assign T1078 = T1071[4'he:4'he];
  assign T1079 = T1071[5'h1e:4'hf];
  assign T1080 = T1094 ? T1091 : T1081;
  assign T1081 = T1087 ? 1'h0 : T1082;
  assign T1082 = T1083 & T1021;
  assign T1083 = T1085 & T1084;
  assign T1084 = VCRouterStateManagement_4_io_currentState == 3'h4;
  assign T1085 = T1040 | T1086;
  assign T1086 = VCRouterStateManagement_4_io_currentState == 3'h4;
  assign T1087 = T1089 & T1088;
  assign T1088 = ~ RouterRegFile_4_io_readValid;
  assign T1089 = T1090 == 1'h1;
  assign T1090 = RouterBuffer_4_io_deq_bits_x[1'h0:1'h0];
  assign T1091 = T1092 & T1021;
  assign T1092 = T1085 & T1093;
  assign T1093 = 3'h3 <= VCRouterStateManagement_4_io_currentState;
  assign T1094 = T1098 & T1095;
  assign T1095 = T1096 & RouterRegFile_4_io_readValid;
  assign T1096 = T1097 == 1'h1;
  assign T1097 = RouterBuffer_4_io_deq_bits_x[1'h0:1'h0];
  assign T1098 = T1087 ^ 1'h1;
  assign T1099 = io_inChannels_2_flitValid & T114;
  assign T1100 = T1101 & RouterRegFile_4_io_readValid;
  assign T1101 = RouterRegFile_4_io_rvPipelineReg_0 ^ 1'h1;
  assign T1102 = T1104 & T1103;
  assign T1103 = VCRouterStateManagement_4_io_currentState == 3'h2;
  assign T1104 = RouterRegFile_4_io_rvPipelineReg_0 & vcAllocator_io_resources_4_valid;
  assign T1105 = T1107 & T1106;
  assign T1106 = VCRouterStateManagement_4_io_currentState == 3'h3;
  assign T1107 = RouterRegFile_4_io_rvPipelineReg_1 & T1040;
  assign T3153 = {24'h0, T1108};
  assign T1108 = T1109;
  assign T1109 = {T1113, T1110};
  assign T1110 = {T1112, T1111};
  assign T1111 = {CMeshDOR_4_io_outHeadFlit_destination_0, CMeshDOR_4_io_outHeadFlit_priorityLevel};
  assign T1112 = {CMeshDOR_4_io_outHeadFlit_destination_2, CMeshDOR_4_io_outHeadFlit_destination_1};
  assign T1113 = {T1115, T1114};
  assign T1114 = {CMeshDOR_4_io_outHeadFlit_vcPort, CMeshDOR_4_io_outHeadFlit_packetType};
  assign T1115 = {CMeshDOR_4_io_outHeadFlit_packetID, CMeshDOR_4_io_outHeadFlit_isTail};
  assign T1116 = T1118 & T1117;
  assign T1117 = VCRouterStateManagement_4_io_currentState == 3'h4;
  assign T1118 = T1119 & T1021;
  assign T1119 = T1085 & flitsAreTail_4;
  assign flitsAreTail_4 = T1120;
  assign T1120 = T1121 & RouterBuffer_4_io_deq_valid;
  assign T1121 = T1122;
  assign T1122 = T1127 ? T1125 : T1123;
  assign T1123 = T1124[6'h25:6'h25];
  assign T1124 = RouterBuffer_4_io_deq_bits_x[6'h36:1'h1];
  assign T1125 = T1126[4'he:4'he];
  assign T1126 = RouterBuffer_4_io_deq_bits_x[5'h1f:1'h1];
  assign T1127 = T1128 == 1'h1;
  assign T1128 = RouterBuffer_4_io_deq_bits_x[1'h0:1'h0];
  assign T1129 = T1130 ? T1099 : 1'h0;
  assign T1130 = T1131 == 1'h1;
  assign T1131 = io_inChannels_2_flit_x[1'h0:1'h0];
  assign T1132 = T1130 ? T1133 : 55'h0;
  assign T1133 = io_inChannels_2_flit_x;
  assign T1134 = T1094 ? T1140 : T1135;
  assign T1135 = T1087 ? 1'h0 : T1136;
  assign T1136 = T1137 & RouterBuffer_4_io_deq_valid;
  assign T1137 = T1138 & T1021;
  assign T1138 = T1085 & T1139;
  assign T1139 = VCRouterStateManagement_4_io_currentState == 3'h4;
  assign T1140 = T1141 & RouterBuffer_4_io_deq_valid;
  assign T1141 = T1142 & T1021;
  assign T1142 = T1085 & T1143;
  assign T1143 = 3'h3 <= VCRouterStateManagement_4_io_currentState;
  assign T1144 = T1145;
  assign T1145 = io_inChannels_1_flit_x;
  assign T3154 = R1146[1'h0:1'h0];
  assign T3155 = reset ? 55'h0 : T1147;
  assign T1147 = T1148 ? T3156 : R1146;
  assign T3156 = {51'h0, vcAllocator_io_chosens_3};
  assign T1148 = T1149 & vcAllocator_io_resources_3_valid;
  assign T1149 = VCRouterStateManagement_3_io_currentState == 3'h2;
  assign T1150 = T1151;
  assign T1151 = RouterBuffer_3_io_deq_bits_x;
  assign T1152 = T1164 | T1153;
  assign T1153 = T1154 == 2'h1;
  assign T1154 = T1163 ? VCRouterOutputStateManagement_4_io_currentState : T1155;
  assign T1155 = T1162 ? T1160 : T1156;
  assign T1156 = T1157 ? VCRouterOutputStateManagement_1_io_currentState : VCRouterOutputStateManagement_io_currentState;
  assign T1157 = T1158[1'h0:1'h0];
  assign T1158 = R1159;
  assign T3157 = reset ? 3'h0 : CMeshDOR_3_io_result;
  assign T1160 = T1161 ? VCRouterOutputStateManagement_3_io_currentState : VCRouterOutputStateManagement_2_io_currentState;
  assign T1161 = T1158[1'h0:1'h0];
  assign T1162 = T1158[1'h1:1'h1];
  assign T1163 = T1158[2'h2:2'h2];
  assign T1164 = T1154 == 2'h2;
  assign T1165 = T1183 ? T1175 : T1166;
  assign T1166 = T1174 ? creditConsReady_4_0 : T1167;
  assign T1167 = T1173 ? T1171 : T1168;
  assign T1168 = T1169 ? creditConsReady_1_0 : creditConsReady_0_0;
  assign T1169 = T1170[1'h0:1'h0];
  assign T1170 = R1159;
  assign T1171 = T1172 ? creditConsReady_3_0 : creditConsReady_2_0;
  assign T1172 = T1170[1'h0:1'h0];
  assign T1173 = T1170[1'h1:1'h1];
  assign T1174 = T1170[2'h2:2'h2];
  assign T1175 = T1182 ? creditConsReady_4_1 : T1176;
  assign T1176 = T1181 ? T1179 : T1177;
  assign T1177 = T1178 ? creditConsReady_1_1 : creditConsReady_0_1;
  assign T1178 = T1170[1'h0:1'h0];
  assign T1179 = T1180 ? creditConsReady_3_1 : creditConsReady_2_1;
  assign T1180 = T1170[1'h0:1'h0];
  assign T1181 = T1170[1'h1:1'h1];
  assign T1182 = T1170[2'h2:2'h2];
  assign T1183 = T3158;
  assign T3158 = R1146[1'h0:1'h0];
  assign T1184 = T1195 & T1185;
  assign T1185 = T1186 == 4'h3;
  assign T1186 = T1194 ? swAllocator_io_chosens_4 : T1187;
  assign T1187 = T1193 ? T1191 : T1188;
  assign T1188 = T1189 ? swAllocator_io_chosens_1 : swAllocator_io_chosens_0;
  assign T1189 = T1190[1'h0:1'h0];
  assign T1190 = R1159;
  assign T1191 = T1192 ? swAllocator_io_chosens_3 : swAllocator_io_chosens_2;
  assign T1192 = T1190[1'h0:1'h0];
  assign T1193 = T1190[1'h1:1'h1];
  assign T1194 = T1190[2'h2:2'h2];
  assign T1195 = T1203 ? swAllocator_io_requests_4_3_grant : T1196;
  assign T1196 = T1202 ? T1200 : T1197;
  assign T1197 = T1198 ? swAllocator_io_requests_1_3_grant : swAllocator_io_requests_0_3_grant;
  assign T1198 = T1199[1'h0:1'h0];
  assign T1199 = R1159;
  assign T1200 = T1201 ? swAllocator_io_requests_3_3_grant : swAllocator_io_requests_2_3_grant;
  assign T1201 = T1199[1'h0:1'h0];
  assign T1202 = T1199[1'h1:1'h1];
  assign T1203 = T1199[2'h2:2'h2];
  assign T1204 = RouterBuffer_3_io_deq_valid & T1205;
  assign T1205 = T1206;
  assign T1206 = T1211 ? T1209 : T1207;
  assign T1207 = T1208[6'h25:6'h25];
  assign T1208 = RouterBuffer_3_io_deq_bits_x[6'h36:1'h1];
  assign T1209 = T1210[4'he:4'he];
  assign T1210 = RouterBuffer_3_io_deq_bits_x[5'h1f:1'h1];
  assign T1211 = T1212 == 1'h1;
  assign T1212 = RouterBuffer_3_io_deq_bits_x[1'h0:1'h0];
  assign T3159 = reset ? 1'h0 : RouterBuffer_3_io_deq_valid;
  assign T1214 = T1215[2'h2:1'h0];
  assign T1215 = T1216[5'h1f:1'h1];
  assign T1216 = RouterRegFile_3_io_readData;
  assign T1217 = T1215[3'h4:2'h3];
  assign T1218 = T1215[3'h6:3'h5];
  assign T1219 = T1215[4'h8:3'h7];
  assign T1220 = T1215[4'hc:4'h9];
  assign T1221 = T1215[4'hd:4'hd];
  assign T1222 = T1215[4'he:4'he];
  assign T1223 = T1215[5'h1e:4'hf];
  assign T1224 = T1238 ? T1235 : T1225;
  assign T1225 = T1231 ? 1'h0 : T1226;
  assign T1226 = T1227 & T1165;
  assign T1227 = T1229 & T1228;
  assign T1228 = VCRouterStateManagement_3_io_currentState == 3'h4;
  assign T1229 = T1184 | T1230;
  assign T1230 = VCRouterStateManagement_3_io_currentState == 3'h4;
  assign T1231 = T1233 & T1232;
  assign T1232 = ~ RouterRegFile_3_io_readValid;
  assign T1233 = T1234 == 1'h1;
  assign T1234 = RouterBuffer_3_io_deq_bits_x[1'h0:1'h0];
  assign T1235 = T1236 & T1165;
  assign T1236 = T1229 & T1237;
  assign T1237 = 3'h3 <= VCRouterStateManagement_3_io_currentState;
  assign T1238 = T1242 & T1239;
  assign T1239 = T1240 & RouterRegFile_3_io_readValid;
  assign T1240 = T1241 == 1'h1;
  assign T1241 = RouterBuffer_3_io_deq_bits_x[1'h0:1'h0];
  assign T1242 = T1231 ^ 1'h1;
  assign T1243 = io_inChannels_1_flitValid & T136;
  assign T1244 = T1245 & RouterRegFile_3_io_readValid;
  assign T1245 = RouterRegFile_3_io_rvPipelineReg_0 ^ 1'h1;
  assign T1246 = T1248 & T1247;
  assign T1247 = VCRouterStateManagement_3_io_currentState == 3'h2;
  assign T1248 = RouterRegFile_3_io_rvPipelineReg_0 & vcAllocator_io_resources_3_valid;
  assign T1249 = T1251 & T1250;
  assign T1250 = VCRouterStateManagement_3_io_currentState == 3'h3;
  assign T1251 = RouterRegFile_3_io_rvPipelineReg_1 & T1184;
  assign T3160 = {24'h0, T1252};
  assign T1252 = T1253;
  assign T1253 = {T1257, T1254};
  assign T1254 = {T1256, T1255};
  assign T1255 = {CMeshDOR_3_io_outHeadFlit_destination_0, CMeshDOR_3_io_outHeadFlit_priorityLevel};
  assign T1256 = {CMeshDOR_3_io_outHeadFlit_destination_2, CMeshDOR_3_io_outHeadFlit_destination_1};
  assign T1257 = {T1259, T1258};
  assign T1258 = {CMeshDOR_3_io_outHeadFlit_vcPort, CMeshDOR_3_io_outHeadFlit_packetType};
  assign T1259 = {CMeshDOR_3_io_outHeadFlit_packetID, CMeshDOR_3_io_outHeadFlit_isTail};
  assign T1260 = T1262 & T1261;
  assign T1261 = VCRouterStateManagement_3_io_currentState == 3'h4;
  assign T1262 = T1263 & T1165;
  assign T1263 = T1229 & flitsAreTail_3;
  assign flitsAreTail_3 = T1264;
  assign T1264 = T1265 & RouterBuffer_3_io_deq_valid;
  assign T1265 = T1266;
  assign T1266 = T1271 ? T1269 : T1267;
  assign T1267 = T1268[6'h25:6'h25];
  assign T1268 = RouterBuffer_3_io_deq_bits_x[6'h36:1'h1];
  assign T1269 = T1270[4'he:4'he];
  assign T1270 = RouterBuffer_3_io_deq_bits_x[5'h1f:1'h1];
  assign T1271 = T1272 == 1'h1;
  assign T1272 = RouterBuffer_3_io_deq_bits_x[1'h0:1'h0];
  assign T1273 = T1274 ? T1243 : 1'h0;
  assign T1274 = T1275 == 1'h1;
  assign T1275 = io_inChannels_1_flit_x[1'h0:1'h0];
  assign T1276 = T1274 ? T1277 : 55'h0;
  assign T1277 = io_inChannels_1_flit_x;
  assign T1278 = T1238 ? T1284 : T1279;
  assign T1279 = T1231 ? 1'h0 : T1280;
  assign T1280 = T1281 & RouterBuffer_3_io_deq_valid;
  assign T1281 = T1282 & T1165;
  assign T1282 = T1229 & T1283;
  assign T1283 = VCRouterStateManagement_3_io_currentState == 3'h4;
  assign T1284 = T1285 & RouterBuffer_3_io_deq_valid;
  assign T1285 = T1286 & T1165;
  assign T1286 = T1229 & T1287;
  assign T1287 = 3'h3 <= VCRouterStateManagement_3_io_currentState;
  assign T1288 = T1289;
  assign T1289 = io_inChannels_1_flit_x;
  assign T3161 = R1290[1'h0:1'h0];
  assign T3162 = reset ? 55'h0 : T1291;
  assign T1291 = T1292 ? T3163 : R1290;
  assign T3163 = {51'h0, vcAllocator_io_chosens_2};
  assign T1292 = T1293 & vcAllocator_io_resources_2_valid;
  assign T1293 = VCRouterStateManagement_2_io_currentState == 3'h2;
  assign T1294 = T1295;
  assign T1295 = RouterBuffer_2_io_deq_bits_x;
  assign T1296 = T1308 | T1297;
  assign T1297 = T1298 == 2'h1;
  assign T1298 = T1307 ? VCRouterOutputStateManagement_4_io_currentState : T1299;
  assign T1299 = T1306 ? T1304 : T1300;
  assign T1300 = T1301 ? VCRouterOutputStateManagement_1_io_currentState : VCRouterOutputStateManagement_io_currentState;
  assign T1301 = T1302[1'h0:1'h0];
  assign T1302 = R1303;
  assign T3164 = reset ? 3'h0 : CMeshDOR_2_io_result;
  assign T1304 = T1305 ? VCRouterOutputStateManagement_3_io_currentState : VCRouterOutputStateManagement_2_io_currentState;
  assign T1305 = T1302[1'h0:1'h0];
  assign T1306 = T1302[1'h1:1'h1];
  assign T1307 = T1302[2'h2:2'h2];
  assign T1308 = T1298 == 2'h2;
  assign T1309 = T1327 ? T1319 : T1310;
  assign T1310 = T1318 ? creditConsReady_4_0 : T1311;
  assign T1311 = T1317 ? T1315 : T1312;
  assign T1312 = T1313 ? creditConsReady_1_0 : creditConsReady_0_0;
  assign T1313 = T1314[1'h0:1'h0];
  assign T1314 = R1303;
  assign T1315 = T1316 ? creditConsReady_3_0 : creditConsReady_2_0;
  assign T1316 = T1314[1'h0:1'h0];
  assign T1317 = T1314[1'h1:1'h1];
  assign T1318 = T1314[2'h2:2'h2];
  assign T1319 = T1326 ? creditConsReady_4_1 : T1320;
  assign T1320 = T1325 ? T1323 : T1321;
  assign T1321 = T1322 ? creditConsReady_1_1 : creditConsReady_0_1;
  assign T1322 = T1314[1'h0:1'h0];
  assign T1323 = T1324 ? creditConsReady_3_1 : creditConsReady_2_1;
  assign T1324 = T1314[1'h0:1'h0];
  assign T1325 = T1314[1'h1:1'h1];
  assign T1326 = T1314[2'h2:2'h2];
  assign T1327 = T3165;
  assign T3165 = R1290[1'h0:1'h0];
  assign T1328 = T1339 & T1329;
  assign T1329 = T1330 == 4'h2;
  assign T1330 = T1338 ? swAllocator_io_chosens_4 : T1331;
  assign T1331 = T1337 ? T1335 : T1332;
  assign T1332 = T1333 ? swAllocator_io_chosens_1 : swAllocator_io_chosens_0;
  assign T1333 = T1334[1'h0:1'h0];
  assign T1334 = R1303;
  assign T1335 = T1336 ? swAllocator_io_chosens_3 : swAllocator_io_chosens_2;
  assign T1336 = T1334[1'h0:1'h0];
  assign T1337 = T1334[1'h1:1'h1];
  assign T1338 = T1334[2'h2:2'h2];
  assign T1339 = T1347 ? swAllocator_io_requests_4_2_grant : T1340;
  assign T1340 = T1346 ? T1344 : T1341;
  assign T1341 = T1342 ? swAllocator_io_requests_1_2_grant : swAllocator_io_requests_0_2_grant;
  assign T1342 = T1343[1'h0:1'h0];
  assign T1343 = R1303;
  assign T1344 = T1345 ? swAllocator_io_requests_3_2_grant : swAllocator_io_requests_2_2_grant;
  assign T1345 = T1343[1'h0:1'h0];
  assign T1346 = T1343[1'h1:1'h1];
  assign T1347 = T1343[2'h2:2'h2];
  assign T1348 = RouterBuffer_2_io_deq_valid & T1349;
  assign T1349 = T1350;
  assign T1350 = T1355 ? T1353 : T1351;
  assign T1351 = T1352[6'h25:6'h25];
  assign T1352 = RouterBuffer_2_io_deq_bits_x[6'h36:1'h1];
  assign T1353 = T1354[4'he:4'he];
  assign T1354 = RouterBuffer_2_io_deq_bits_x[5'h1f:1'h1];
  assign T1355 = T1356 == 1'h1;
  assign T1356 = RouterBuffer_2_io_deq_bits_x[1'h0:1'h0];
  assign T3166 = reset ? 1'h0 : RouterBuffer_2_io_deq_valid;
  assign T1358 = T1359[2'h2:1'h0];
  assign T1359 = T1360[5'h1f:1'h1];
  assign T1360 = RouterRegFile_2_io_readData;
  assign T1361 = T1359[3'h4:2'h3];
  assign T1362 = T1359[3'h6:3'h5];
  assign T1363 = T1359[4'h8:3'h7];
  assign T1364 = T1359[4'hc:4'h9];
  assign T1365 = T1359[4'hd:4'hd];
  assign T1366 = T1359[4'he:4'he];
  assign T1367 = T1359[5'h1e:4'hf];
  assign T1368 = T1382 ? T1379 : T1369;
  assign T1369 = T1375 ? 1'h0 : T1370;
  assign T1370 = T1371 & T1309;
  assign T1371 = T1373 & T1372;
  assign T1372 = VCRouterStateManagement_2_io_currentState == 3'h4;
  assign T1373 = T1328 | T1374;
  assign T1374 = VCRouterStateManagement_2_io_currentState == 3'h4;
  assign T1375 = T1377 & T1376;
  assign T1376 = ~ RouterRegFile_2_io_readValid;
  assign T1377 = T1378 == 1'h1;
  assign T1378 = RouterBuffer_2_io_deq_bits_x[1'h0:1'h0];
  assign T1379 = T1380 & T1309;
  assign T1380 = T1373 & T1381;
  assign T1381 = 3'h3 <= VCRouterStateManagement_2_io_currentState;
  assign T1382 = T1386 & T1383;
  assign T1383 = T1384 & RouterRegFile_2_io_readValid;
  assign T1384 = T1385 == 1'h1;
  assign T1385 = RouterBuffer_2_io_deq_bits_x[1'h0:1'h0];
  assign T1386 = T1375 ^ 1'h1;
  assign T1387 = io_inChannels_1_flitValid & T158;
  assign T1388 = T1389 & RouterRegFile_2_io_readValid;
  assign T1389 = RouterRegFile_2_io_rvPipelineReg_0 ^ 1'h1;
  assign T1390 = T1392 & T1391;
  assign T1391 = VCRouterStateManagement_2_io_currentState == 3'h2;
  assign T1392 = RouterRegFile_2_io_rvPipelineReg_0 & vcAllocator_io_resources_2_valid;
  assign T1393 = T1395 & T1394;
  assign T1394 = VCRouterStateManagement_2_io_currentState == 3'h3;
  assign T1395 = RouterRegFile_2_io_rvPipelineReg_1 & T1328;
  assign T3167 = {24'h0, T1396};
  assign T1396 = T1397;
  assign T1397 = {T1401, T1398};
  assign T1398 = {T1400, T1399};
  assign T1399 = {CMeshDOR_2_io_outHeadFlit_destination_0, CMeshDOR_2_io_outHeadFlit_priorityLevel};
  assign T1400 = {CMeshDOR_2_io_outHeadFlit_destination_2, CMeshDOR_2_io_outHeadFlit_destination_1};
  assign T1401 = {T1403, T1402};
  assign T1402 = {CMeshDOR_2_io_outHeadFlit_vcPort, CMeshDOR_2_io_outHeadFlit_packetType};
  assign T1403 = {CMeshDOR_2_io_outHeadFlit_packetID, CMeshDOR_2_io_outHeadFlit_isTail};
  assign T1404 = T1406 & T1405;
  assign T1405 = VCRouterStateManagement_2_io_currentState == 3'h4;
  assign T1406 = T1407 & T1309;
  assign T1407 = T1373 & flitsAreTail_2;
  assign flitsAreTail_2 = T1408;
  assign T1408 = T1409 & RouterBuffer_2_io_deq_valid;
  assign T1409 = T1410;
  assign T1410 = T1415 ? T1413 : T1411;
  assign T1411 = T1412[6'h25:6'h25];
  assign T1412 = RouterBuffer_2_io_deq_bits_x[6'h36:1'h1];
  assign T1413 = T1414[4'he:4'he];
  assign T1414 = RouterBuffer_2_io_deq_bits_x[5'h1f:1'h1];
  assign T1415 = T1416 == 1'h1;
  assign T1416 = RouterBuffer_2_io_deq_bits_x[1'h0:1'h0];
  assign T1417 = T1418 ? T1387 : 1'h0;
  assign T1418 = T1419 == 1'h1;
  assign T1419 = io_inChannels_1_flit_x[1'h0:1'h0];
  assign T1420 = T1418 ? T1421 : 55'h0;
  assign T1421 = io_inChannels_1_flit_x;
  assign T1422 = T1382 ? T1428 : T1423;
  assign T1423 = T1375 ? 1'h0 : T1424;
  assign T1424 = T1425 & RouterBuffer_2_io_deq_valid;
  assign T1425 = T1426 & T1309;
  assign T1426 = T1373 & T1427;
  assign T1427 = VCRouterStateManagement_2_io_currentState == 3'h4;
  assign T1428 = T1429 & RouterBuffer_2_io_deq_valid;
  assign T1429 = T1430 & T1309;
  assign T1430 = T1373 & T1431;
  assign T1431 = 3'h3 <= VCRouterStateManagement_2_io_currentState;
  assign T1432 = T1433;
  assign T1433 = io_inChannels_0_flit_x;
  assign T3168 = R1434[1'h0:1'h0];
  assign T3169 = reset ? 55'h0 : T1435;
  assign T1435 = T1436 ? T3170 : R1434;
  assign T3170 = {51'h0, vcAllocator_io_chosens_1};
  assign T1436 = T1437 & vcAllocator_io_resources_1_valid;
  assign T1437 = VCRouterStateManagement_1_io_currentState == 3'h2;
  assign T1438 = T1439;
  assign T1439 = RouterBuffer_1_io_deq_bits_x;
  assign T1440 = T1452 | T1441;
  assign T1441 = T1442 == 2'h1;
  assign T1442 = T1451 ? VCRouterOutputStateManagement_4_io_currentState : T1443;
  assign T1443 = T1450 ? T1448 : T1444;
  assign T1444 = T1445 ? VCRouterOutputStateManagement_1_io_currentState : VCRouterOutputStateManagement_io_currentState;
  assign T1445 = T1446[1'h0:1'h0];
  assign T1446 = R1447;
  assign T3171 = reset ? 3'h0 : CMeshDOR_1_io_result;
  assign T1448 = T1449 ? VCRouterOutputStateManagement_3_io_currentState : VCRouterOutputStateManagement_2_io_currentState;
  assign T1449 = T1446[1'h0:1'h0];
  assign T1450 = T1446[1'h1:1'h1];
  assign T1451 = T1446[2'h2:2'h2];
  assign T1452 = T1442 == 2'h2;
  assign T1453 = T1471 ? T1463 : T1454;
  assign T1454 = T1462 ? creditConsReady_4_0 : T1455;
  assign T1455 = T1461 ? T1459 : T1456;
  assign T1456 = T1457 ? creditConsReady_1_0 : creditConsReady_0_0;
  assign T1457 = T1458[1'h0:1'h0];
  assign T1458 = R1447;
  assign T1459 = T1460 ? creditConsReady_3_0 : creditConsReady_2_0;
  assign T1460 = T1458[1'h0:1'h0];
  assign T1461 = T1458[1'h1:1'h1];
  assign T1462 = T1458[2'h2:2'h2];
  assign T1463 = T1470 ? creditConsReady_4_1 : T1464;
  assign T1464 = T1469 ? T1467 : T1465;
  assign T1465 = T1466 ? creditConsReady_1_1 : creditConsReady_0_1;
  assign T1466 = T1458[1'h0:1'h0];
  assign T1467 = T1468 ? creditConsReady_3_1 : creditConsReady_2_1;
  assign T1468 = T1458[1'h0:1'h0];
  assign T1469 = T1458[1'h1:1'h1];
  assign T1470 = T1458[2'h2:2'h2];
  assign T1471 = T3172;
  assign T3172 = R1434[1'h0:1'h0];
  assign T1472 = T1483 & T1473;
  assign T1473 = T1474 == 4'h1;
  assign T1474 = T1482 ? swAllocator_io_chosens_4 : T1475;
  assign T1475 = T1481 ? T1479 : T1476;
  assign T1476 = T1477 ? swAllocator_io_chosens_1 : swAllocator_io_chosens_0;
  assign T1477 = T1478[1'h0:1'h0];
  assign T1478 = R1447;
  assign T1479 = T1480 ? swAllocator_io_chosens_3 : swAllocator_io_chosens_2;
  assign T1480 = T1478[1'h0:1'h0];
  assign T1481 = T1478[1'h1:1'h1];
  assign T1482 = T1478[2'h2:2'h2];
  assign T1483 = T1491 ? swAllocator_io_requests_4_1_grant : T1484;
  assign T1484 = T1490 ? T1488 : T1485;
  assign T1485 = T1486 ? swAllocator_io_requests_1_1_grant : swAllocator_io_requests_0_1_grant;
  assign T1486 = T1487[1'h0:1'h0];
  assign T1487 = R1447;
  assign T1488 = T1489 ? swAllocator_io_requests_3_1_grant : swAllocator_io_requests_2_1_grant;
  assign T1489 = T1487[1'h0:1'h0];
  assign T1490 = T1487[1'h1:1'h1];
  assign T1491 = T1487[2'h2:2'h2];
  assign T1492 = RouterBuffer_1_io_deq_valid & T1493;
  assign T1493 = T1494;
  assign T1494 = T1499 ? T1497 : T1495;
  assign T1495 = T1496[6'h25:6'h25];
  assign T1496 = RouterBuffer_1_io_deq_bits_x[6'h36:1'h1];
  assign T1497 = T1498[4'he:4'he];
  assign T1498 = RouterBuffer_1_io_deq_bits_x[5'h1f:1'h1];
  assign T1499 = T1500 == 1'h1;
  assign T1500 = RouterBuffer_1_io_deq_bits_x[1'h0:1'h0];
  assign T3173 = reset ? 1'h0 : RouterBuffer_1_io_deq_valid;
  assign T1502 = T1503[2'h2:1'h0];
  assign T1503 = T1504[5'h1f:1'h1];
  assign T1504 = RouterRegFile_1_io_readData;
  assign T1505 = T1503[3'h4:2'h3];
  assign T1506 = T1503[3'h6:3'h5];
  assign T1507 = T1503[4'h8:3'h7];
  assign T1508 = T1503[4'hc:4'h9];
  assign T1509 = T1503[4'hd:4'hd];
  assign T1510 = T1503[4'he:4'he];
  assign T1511 = T1503[5'h1e:4'hf];
  assign T1512 = T1526 ? T1523 : T1513;
  assign T1513 = T1519 ? 1'h0 : T1514;
  assign T1514 = T1515 & T1453;
  assign T1515 = T1517 & T1516;
  assign T1516 = VCRouterStateManagement_1_io_currentState == 3'h4;
  assign T1517 = T1472 | T1518;
  assign T1518 = VCRouterStateManagement_1_io_currentState == 3'h4;
  assign T1519 = T1521 & T1520;
  assign T1520 = ~ RouterRegFile_1_io_readValid;
  assign T1521 = T1522 == 1'h1;
  assign T1522 = RouterBuffer_1_io_deq_bits_x[1'h0:1'h0];
  assign T1523 = T1524 & T1453;
  assign T1524 = T1517 & T1525;
  assign T1525 = 3'h3 <= VCRouterStateManagement_1_io_currentState;
  assign T1526 = T1530 & T1527;
  assign T1527 = T1528 & RouterRegFile_1_io_readValid;
  assign T1528 = T1529 == 1'h1;
  assign T1529 = RouterBuffer_1_io_deq_bits_x[1'h0:1'h0];
  assign T1530 = T1519 ^ 1'h1;
  assign T1531 = io_inChannels_0_flitValid & T180;
  assign T1532 = T1533 & RouterRegFile_1_io_readValid;
  assign T1533 = RouterRegFile_1_io_rvPipelineReg_0 ^ 1'h1;
  assign T1534 = T1536 & T1535;
  assign T1535 = VCRouterStateManagement_1_io_currentState == 3'h2;
  assign T1536 = RouterRegFile_1_io_rvPipelineReg_0 & vcAllocator_io_resources_1_valid;
  assign T1537 = T1539 & T1538;
  assign T1538 = VCRouterStateManagement_1_io_currentState == 3'h3;
  assign T1539 = RouterRegFile_1_io_rvPipelineReg_1 & T1472;
  assign T3174 = {24'h0, T1540};
  assign T1540 = T1541;
  assign T1541 = {T1545, T1542};
  assign T1542 = {T1544, T1543};
  assign T1543 = {CMeshDOR_1_io_outHeadFlit_destination_0, CMeshDOR_1_io_outHeadFlit_priorityLevel};
  assign T1544 = {CMeshDOR_1_io_outHeadFlit_destination_2, CMeshDOR_1_io_outHeadFlit_destination_1};
  assign T1545 = {T1547, T1546};
  assign T1546 = {CMeshDOR_1_io_outHeadFlit_vcPort, CMeshDOR_1_io_outHeadFlit_packetType};
  assign T1547 = {CMeshDOR_1_io_outHeadFlit_packetID, CMeshDOR_1_io_outHeadFlit_isTail};
  assign T1548 = T1550 & T1549;
  assign T1549 = VCRouterStateManagement_1_io_currentState == 3'h4;
  assign T1550 = T1551 & T1453;
  assign T1551 = T1517 & flitsAreTail_1;
  assign flitsAreTail_1 = T1552;
  assign T1552 = T1553 & RouterBuffer_1_io_deq_valid;
  assign T1553 = T1554;
  assign T1554 = T1559 ? T1557 : T1555;
  assign T1555 = T1556[6'h25:6'h25];
  assign T1556 = RouterBuffer_1_io_deq_bits_x[6'h36:1'h1];
  assign T1557 = T1558[4'he:4'he];
  assign T1558 = RouterBuffer_1_io_deq_bits_x[5'h1f:1'h1];
  assign T1559 = T1560 == 1'h1;
  assign T1560 = RouterBuffer_1_io_deq_bits_x[1'h0:1'h0];
  assign T1561 = T1562 ? T1531 : 1'h0;
  assign T1562 = T1563 == 1'h1;
  assign T1563 = io_inChannels_0_flit_x[1'h0:1'h0];
  assign T1564 = T1562 ? T1565 : 55'h0;
  assign T1565 = io_inChannels_0_flit_x;
  assign T1566 = T1526 ? T1572 : T1567;
  assign T1567 = T1519 ? 1'h0 : T1568;
  assign T1568 = T1569 & RouterBuffer_1_io_deq_valid;
  assign T1569 = T1570 & T1453;
  assign T1570 = T1517 & T1571;
  assign T1571 = VCRouterStateManagement_1_io_currentState == 3'h4;
  assign T1572 = T1573 & RouterBuffer_1_io_deq_valid;
  assign T1573 = T1574 & T1453;
  assign T1574 = T1517 & T1575;
  assign T1575 = 3'h3 <= VCRouterStateManagement_1_io_currentState;
  assign T1576 = T1577;
  assign T1577 = io_inChannels_0_flit_x;
  assign T3175 = R1578[1'h0:1'h0];
  assign T3176 = reset ? 55'h0 : T1579;
  assign T1579 = T1580 ? T3177 : R1578;
  assign T3177 = {51'h0, vcAllocator_io_chosens_0};
  assign T1580 = T1581 & vcAllocator_io_resources_0_valid;
  assign T1581 = VCRouterStateManagement_io_currentState == 3'h2;
  assign T1582 = T1583;
  assign T1583 = RouterBuffer_io_deq_bits_x;
  assign T1584 = T1596 | T1585;
  assign T1585 = T1586 == 2'h1;
  assign T1586 = T1595 ? VCRouterOutputStateManagement_4_io_currentState : T1587;
  assign T1587 = T1594 ? T1592 : T1588;
  assign T1588 = T1589 ? VCRouterOutputStateManagement_1_io_currentState : VCRouterOutputStateManagement_io_currentState;
  assign T1589 = T1590[1'h0:1'h0];
  assign T1590 = R1591;
  assign T3178 = reset ? 3'h0 : CMeshDOR_io_result;
  assign T1592 = T1593 ? VCRouterOutputStateManagement_3_io_currentState : VCRouterOutputStateManagement_2_io_currentState;
  assign T1593 = T1590[1'h0:1'h0];
  assign T1594 = T1590[1'h1:1'h1];
  assign T1595 = T1590[2'h2:2'h2];
  assign T1596 = T1586 == 2'h2;
  assign T1597 = T1615 ? T1607 : T1598;
  assign T1598 = T1606 ? creditConsReady_4_0 : T1599;
  assign T1599 = T1605 ? T1603 : T1600;
  assign T1600 = T1601 ? creditConsReady_1_0 : creditConsReady_0_0;
  assign T1601 = T1602[1'h0:1'h0];
  assign T1602 = R1591;
  assign T1603 = T1604 ? creditConsReady_3_0 : creditConsReady_2_0;
  assign T1604 = T1602[1'h0:1'h0];
  assign T1605 = T1602[1'h1:1'h1];
  assign T1606 = T1602[2'h2:2'h2];
  assign T1607 = T1614 ? creditConsReady_4_1 : T1608;
  assign T1608 = T1613 ? T1611 : T1609;
  assign T1609 = T1610 ? creditConsReady_1_1 : creditConsReady_0_1;
  assign T1610 = T1602[1'h0:1'h0];
  assign T1611 = T1612 ? creditConsReady_3_1 : creditConsReady_2_1;
  assign T1612 = T1602[1'h0:1'h0];
  assign T1613 = T1602[1'h1:1'h1];
  assign T1614 = T1602[2'h2:2'h2];
  assign T1615 = T3179;
  assign T3179 = R1578[1'h0:1'h0];
  assign T1616 = T1627 & T1617;
  assign T1617 = T1618 == 4'h0;
  assign T1618 = T1626 ? swAllocator_io_chosens_4 : T1619;
  assign T1619 = T1625 ? T1623 : T1620;
  assign T1620 = T1621 ? swAllocator_io_chosens_1 : swAllocator_io_chosens_0;
  assign T1621 = T1622[1'h0:1'h0];
  assign T1622 = R1591;
  assign T1623 = T1624 ? swAllocator_io_chosens_3 : swAllocator_io_chosens_2;
  assign T1624 = T1622[1'h0:1'h0];
  assign T1625 = T1622[1'h1:1'h1];
  assign T1626 = T1622[2'h2:2'h2];
  assign T1627 = T1635 ? swAllocator_io_requests_4_0_grant : T1628;
  assign T1628 = T1634 ? T1632 : T1629;
  assign T1629 = T1630 ? swAllocator_io_requests_1_0_grant : swAllocator_io_requests_0_0_grant;
  assign T1630 = T1631[1'h0:1'h0];
  assign T1631 = R1591;
  assign T1632 = T1633 ? swAllocator_io_requests_3_0_grant : swAllocator_io_requests_2_0_grant;
  assign T1633 = T1631[1'h0:1'h0];
  assign T1634 = T1631[1'h1:1'h1];
  assign T1635 = T1631[2'h2:2'h2];
  assign T1636 = RouterBuffer_io_deq_valid & T1637;
  assign T1637 = T1638;
  assign T1638 = T1643 ? T1641 : T1639;
  assign T1639 = T1640[6'h25:6'h25];
  assign T1640 = RouterBuffer_io_deq_bits_x[6'h36:1'h1];
  assign T1641 = T1642[4'he:4'he];
  assign T1642 = RouterBuffer_io_deq_bits_x[5'h1f:1'h1];
  assign T1643 = T1644 == 1'h1;
  assign T1644 = RouterBuffer_io_deq_bits_x[1'h0:1'h0];
  assign T3180 = reset ? 1'h0 : RouterBuffer_io_deq_valid;
  assign T1646 = T1647[2'h2:1'h0];
  assign T1647 = T1648[5'h1f:1'h1];
  assign T1648 = RouterRegFile_io_readData;
  assign T1649 = T1647[3'h4:2'h3];
  assign T1650 = T1647[3'h6:3'h5];
  assign T1651 = T1647[4'h8:3'h7];
  assign T1652 = T1647[4'hc:4'h9];
  assign T1653 = T1647[4'hd:4'hd];
  assign T1654 = T1647[4'he:4'he];
  assign T1655 = T1647[5'h1e:4'hf];
  assign T1656 = T1670 ? T1667 : T1657;
  assign T1657 = T1663 ? 1'h0 : T1658;
  assign T1658 = T1659 & T1597;
  assign T1659 = T1661 & T1660;
  assign T1660 = VCRouterStateManagement_io_currentState == 3'h4;
  assign T1661 = T1616 | T1662;
  assign T1662 = VCRouterStateManagement_io_currentState == 3'h4;
  assign T1663 = T1665 & T1664;
  assign T1664 = ~ RouterRegFile_io_readValid;
  assign T1665 = T1666 == 1'h1;
  assign T1666 = RouterBuffer_io_deq_bits_x[1'h0:1'h0];
  assign T1667 = T1668 & T1597;
  assign T1668 = T1661 & T1669;
  assign T1669 = 3'h3 <= VCRouterStateManagement_io_currentState;
  assign T1670 = T1674 & T1671;
  assign T1671 = T1672 & RouterRegFile_io_readValid;
  assign T1672 = T1673 == 1'h1;
  assign T1673 = RouterBuffer_io_deq_bits_x[1'h0:1'h0];
  assign T1674 = T1663 ^ 1'h1;
  assign T1675 = io_inChannels_0_flitValid & T202;
  assign T1676 = T1677 & RouterRegFile_io_readValid;
  assign T1677 = RouterRegFile_io_rvPipelineReg_0 ^ 1'h1;
  assign T1678 = T1680 & T1679;
  assign T1679 = VCRouterStateManagement_io_currentState == 3'h2;
  assign T1680 = RouterRegFile_io_rvPipelineReg_0 & vcAllocator_io_resources_0_valid;
  assign T1681 = T1683 & T1682;
  assign T1682 = VCRouterStateManagement_io_currentState == 3'h3;
  assign T1683 = RouterRegFile_io_rvPipelineReg_1 & T1616;
  assign T3181 = {24'h0, T1684};
  assign T1684 = T1685;
  assign T1685 = {T1689, T1686};
  assign T1686 = {T1688, T1687};
  assign T1687 = {CMeshDOR_io_outHeadFlit_destination_0, CMeshDOR_io_outHeadFlit_priorityLevel};
  assign T1688 = {CMeshDOR_io_outHeadFlit_destination_2, CMeshDOR_io_outHeadFlit_destination_1};
  assign T1689 = {T1691, T1690};
  assign T1690 = {CMeshDOR_io_outHeadFlit_vcPort, CMeshDOR_io_outHeadFlit_packetType};
  assign T1691 = {CMeshDOR_io_outHeadFlit_packetID, CMeshDOR_io_outHeadFlit_isTail};
  assign T1692 = T1694 & T1693;
  assign T1693 = VCRouterStateManagement_io_currentState == 3'h4;
  assign T1694 = T1695 & T1597;
  assign T1695 = T1661 & flitsAreTail_0;
  assign flitsAreTail_0 = T1696;
  assign T1696 = T1697 & RouterBuffer_io_deq_valid;
  assign T1697 = T1698;
  assign T1698 = T1703 ? T1701 : T1699;
  assign T1699 = T1700[6'h25:6'h25];
  assign T1700 = RouterBuffer_io_deq_bits_x[6'h36:1'h1];
  assign T1701 = T1702[4'he:4'he];
  assign T1702 = RouterBuffer_io_deq_bits_x[5'h1f:1'h1];
  assign T1703 = T1704 == 1'h1;
  assign T1704 = RouterBuffer_io_deq_bits_x[1'h0:1'h0];
  assign T1705 = T1706 ? T1675 : 1'h0;
  assign T1706 = T1707 == 1'h1;
  assign T1707 = io_inChannels_0_flit_x[1'h0:1'h0];
  assign T1708 = T1706 ? T1709 : 55'h0;
  assign T1709 = io_inChannels_0_flit_x;
  assign T1710 = T1670 ? T1716 : T1711;
  assign T1711 = T1663 ? 1'h0 : T1712;
  assign T1712 = T1713 & RouterBuffer_io_deq_valid;
  assign T1713 = T1714 & T1597;
  assign T1714 = T1661 & T1715;
  assign T1715 = VCRouterStateManagement_io_currentState == 3'h4;
  assign T1716 = T1717 & RouterBuffer_io_deq_valid;
  assign T1717 = T1718 & T1597;
  assign T1718 = T1661 & T1719;
  assign T1719 = 3'h3 <= VCRouterStateManagement_io_currentState;
  assign T1720 = T1721 ? CreditCon_9_io_outCredit : CreditCon_8_io_outCredit;
  assign T1721 = T222;
  assign T1722 = T1723 != 10'h0;
  assign T1723 = T1724;
  assign T1724 = {T1814, T1725};
  assign T1725 = {T1779, T1726};
  assign T1726 = {readyToXmit_2_4, T1727};
  assign T1727 = {readyToXmit_1_4, readyToXmit_0_4};
  assign readyToXmit_0_4 = T1728;
  assign T1728 = T1742 ? T1738 : T1729;
  assign T1729 = T1734 ? T1730 : 1'h0;
  assign T1730 = T1731 & RouterBuffer_io_deq_valid;
  assign T1731 = T1732 & T1597;
  assign T1732 = T1661 & T1733;
  assign T1733 = 3'h3 <= VCRouterStateManagement_io_currentState;
  assign T1734 = T1670 & T1735;
  assign T1735 = T1736[3'h4:3'h4];
  assign T1736 = 1'h1 << T1737;
  assign T1737 = R1591;
  assign T1738 = T1739 & RouterBuffer_io_deq_valid;
  assign T1739 = T1740 & T1597;
  assign T1740 = T1661 & T1741;
  assign T1741 = VCRouterStateManagement_io_currentState == 3'h4;
  assign T1742 = T1743 & T1735;
  assign T1743 = T1744 ^ 1'h1;
  assign T1744 = T1663 | T1671;
  assign readyToXmit_1_4 = T1745;
  assign T1745 = T1759 ? T1755 : T1746;
  assign T1746 = T1751 ? T1747 : 1'h0;
  assign T1747 = T1748 & RouterBuffer_1_io_deq_valid;
  assign T1748 = T1749 & T1453;
  assign T1749 = T1517 & T1750;
  assign T1750 = 3'h3 <= VCRouterStateManagement_1_io_currentState;
  assign T1751 = T1526 & T1752;
  assign T1752 = T1753[3'h4:3'h4];
  assign T1753 = 1'h1 << T1754;
  assign T1754 = R1447;
  assign T1755 = T1756 & RouterBuffer_1_io_deq_valid;
  assign T1756 = T1757 & T1453;
  assign T1757 = T1517 & T1758;
  assign T1758 = VCRouterStateManagement_1_io_currentState == 3'h4;
  assign T1759 = T1760 & T1752;
  assign T1760 = T1761 ^ 1'h1;
  assign T1761 = T1519 | T1527;
  assign readyToXmit_2_4 = T1762;
  assign T1762 = T1776 ? T1772 : T1763;
  assign T1763 = T1768 ? T1764 : 1'h0;
  assign T1764 = T1765 & RouterBuffer_2_io_deq_valid;
  assign T1765 = T1766 & T1309;
  assign T1766 = T1373 & T1767;
  assign T1767 = 3'h3 <= VCRouterStateManagement_2_io_currentState;
  assign T1768 = T1382 & T1769;
  assign T1769 = T1770[3'h4:3'h4];
  assign T1770 = 1'h1 << T1771;
  assign T1771 = R1303;
  assign T1772 = T1773 & RouterBuffer_2_io_deq_valid;
  assign T1773 = T1774 & T1309;
  assign T1774 = T1373 & T1775;
  assign T1775 = VCRouterStateManagement_2_io_currentState == 3'h4;
  assign T1776 = T1777 & T1769;
  assign T1777 = T1778 ^ 1'h1;
  assign T1778 = T1375 | T1383;
  assign T1779 = {readyToXmit_4_4, readyToXmit_3_4};
  assign readyToXmit_3_4 = T1780;
  assign T1780 = T1794 ? T1790 : T1781;
  assign T1781 = T1786 ? T1782 : 1'h0;
  assign T1782 = T1783 & RouterBuffer_3_io_deq_valid;
  assign T1783 = T1784 & T1165;
  assign T1784 = T1229 & T1785;
  assign T1785 = 3'h3 <= VCRouterStateManagement_3_io_currentState;
  assign T1786 = T1238 & T1787;
  assign T1787 = T1788[3'h4:3'h4];
  assign T1788 = 1'h1 << T1789;
  assign T1789 = R1159;
  assign T1790 = T1791 & RouterBuffer_3_io_deq_valid;
  assign T1791 = T1792 & T1165;
  assign T1792 = T1229 & T1793;
  assign T1793 = VCRouterStateManagement_3_io_currentState == 3'h4;
  assign T1794 = T1795 & T1787;
  assign T1795 = T1796 ^ 1'h1;
  assign T1796 = T1231 | T1239;
  assign readyToXmit_4_4 = T1797;
  assign T1797 = T1811 ? T1807 : T1798;
  assign T1798 = T1803 ? T1799 : 1'h0;
  assign T1799 = T1800 & RouterBuffer_4_io_deq_valid;
  assign T1800 = T1801 & T1021;
  assign T1801 = T1085 & T1802;
  assign T1802 = 3'h3 <= VCRouterStateManagement_4_io_currentState;
  assign T1803 = T1094 & T1804;
  assign T1804 = T1805[3'h4:3'h4];
  assign T1805 = 1'h1 << T1806;
  assign T1806 = R1015;
  assign T1807 = T1808 & RouterBuffer_4_io_deq_valid;
  assign T1808 = T1809 & T1021;
  assign T1809 = T1085 & T1810;
  assign T1810 = VCRouterStateManagement_4_io_currentState == 3'h4;
  assign T1811 = T1812 & T1804;
  assign T1812 = T1813 ^ 1'h1;
  assign T1813 = T1087 | T1095;
  assign T1814 = {T1868, T1815};
  assign T1815 = {readyToXmit_7_4, T1816};
  assign T1816 = {readyToXmit_6_4, readyToXmit_5_4};
  assign readyToXmit_5_4 = T1817;
  assign T1817 = T1831 ? T1827 : T1818;
  assign T1818 = T1823 ? T1819 : 1'h0;
  assign T1819 = T1820 & RouterBuffer_5_io_deq_valid;
  assign T1820 = T1821 & T877;
  assign T1821 = T941 & T1822;
  assign T1822 = 3'h3 <= VCRouterStateManagement_5_io_currentState;
  assign T1823 = T950 & T1824;
  assign T1824 = T1825[3'h4:3'h4];
  assign T1825 = 1'h1 << T1826;
  assign T1826 = R871;
  assign T1827 = T1828 & RouterBuffer_5_io_deq_valid;
  assign T1828 = T1829 & T877;
  assign T1829 = T941 & T1830;
  assign T1830 = VCRouterStateManagement_5_io_currentState == 3'h4;
  assign T1831 = T1832 & T1824;
  assign T1832 = T1833 ^ 1'h1;
  assign T1833 = T943 | T951;
  assign readyToXmit_6_4 = T1834;
  assign T1834 = T1848 ? T1844 : T1835;
  assign T1835 = T1840 ? T1836 : 1'h0;
  assign T1836 = T1837 & RouterBuffer_6_io_deq_valid;
  assign T1837 = T1838 & T733;
  assign T1838 = T797 & T1839;
  assign T1839 = 3'h3 <= VCRouterStateManagement_6_io_currentState;
  assign T1840 = T806 & T1841;
  assign T1841 = T1842[3'h4:3'h4];
  assign T1842 = 1'h1 << T1843;
  assign T1843 = R727;
  assign T1844 = T1845 & RouterBuffer_6_io_deq_valid;
  assign T1845 = T1846 & T733;
  assign T1846 = T797 & T1847;
  assign T1847 = VCRouterStateManagement_6_io_currentState == 3'h4;
  assign T1848 = T1849 & T1841;
  assign T1849 = T1850 ^ 1'h1;
  assign T1850 = T799 | T807;
  assign readyToXmit_7_4 = T1851;
  assign T1851 = T1865 ? T1861 : T1852;
  assign T1852 = T1857 ? T1853 : 1'h0;
  assign T1853 = T1854 & RouterBuffer_7_io_deq_valid;
  assign T1854 = T1855 & T589;
  assign T1855 = T653 & T1856;
  assign T1856 = 3'h3 <= VCRouterStateManagement_7_io_currentState;
  assign T1857 = T662 & T1858;
  assign T1858 = T1859[3'h4:3'h4];
  assign T1859 = 1'h1 << T1860;
  assign T1860 = R583;
  assign T1861 = T1862 & RouterBuffer_7_io_deq_valid;
  assign T1862 = T1863 & T589;
  assign T1863 = T653 & T1864;
  assign T1864 = VCRouterStateManagement_7_io_currentState == 3'h4;
  assign T1865 = T1866 & T1858;
  assign T1866 = T1867 ^ 1'h1;
  assign T1867 = T655 | T663;
  assign T1868 = {readyToXmit_9_4, readyToXmit_8_4};
  assign readyToXmit_8_4 = T1869;
  assign T1869 = T1883 ? T1879 : T1870;
  assign T1870 = T1875 ? T1871 : 1'h0;
  assign T1871 = T1872 & RouterBuffer_8_io_deq_valid;
  assign T1872 = T1873 & T445;
  assign T1873 = T509 & T1874;
  assign T1874 = 3'h3 <= VCRouterStateManagement_8_io_currentState;
  assign T1875 = T518 & T1876;
  assign T1876 = T1877[3'h4:3'h4];
  assign T1877 = 1'h1 << T1878;
  assign T1878 = R439;
  assign T1879 = T1880 & RouterBuffer_8_io_deq_valid;
  assign T1880 = T1881 & T445;
  assign T1881 = T509 & T1882;
  assign T1882 = VCRouterStateManagement_8_io_currentState == 3'h4;
  assign T1883 = T1884 & T1876;
  assign T1884 = T1885 ^ 1'h1;
  assign T1885 = T511 | T519;
  assign readyToXmit_9_4 = T1886;
  assign T1886 = T1900 ? T1896 : T1887;
  assign T1887 = T1892 ? T1888 : 1'h0;
  assign T1888 = T1889 & RouterBuffer_9_io_deq_valid;
  assign T1889 = T1890 & T301;
  assign T1890 = T365 & T1891;
  assign T1891 = 3'h3 <= VCRouterStateManagement_9_io_currentState;
  assign T1892 = T374 & T1893;
  assign T1893 = T1894[3'h4:3'h4];
  assign T1894 = 1'h1 << T1895;
  assign T1895 = R295;
  assign T1896 = T1897 & RouterBuffer_9_io_deq_valid;
  assign T1897 = T1898 & T301;
  assign T1898 = T365 & T1899;
  assign T1899 = VCRouterStateManagement_9_io_currentState == 3'h4;
  assign T1900 = T1901 & T1893;
  assign T1901 = T1902 ^ 1'h1;
  assign T1902 = T367 | T375;
  assign T1903 = T1904 ? CreditCon_7_io_outCredit : CreditCon_6_io_outCredit;
  assign T1904 = T234;
  assign T1905 = T1906 != 10'h0;
  assign T1906 = T1907;
  assign T1907 = {T1937, T1908};
  assign T1908 = {T1926, T1909};
  assign T1909 = {readyToXmit_2_3, T1910};
  assign T1910 = {readyToXmit_1_3, readyToXmit_0_3};
  assign readyToXmit_0_3 = T1911;
  assign T1911 = T1915 ? T1738 : T1912;
  assign T1912 = T1913 ? T1730 : 1'h0;
  assign T1913 = T1670 & T1914;
  assign T1914 = T1736[2'h3:2'h3];
  assign T1915 = T1743 & T1914;
  assign readyToXmit_1_3 = T1916;
  assign T1916 = T1920 ? T1755 : T1917;
  assign T1917 = T1918 ? T1747 : 1'h0;
  assign T1918 = T1526 & T1919;
  assign T1919 = T1753[2'h3:2'h3];
  assign T1920 = T1760 & T1919;
  assign readyToXmit_2_3 = T1921;
  assign T1921 = T1925 ? T1772 : T1922;
  assign T1922 = T1923 ? T1764 : 1'h0;
  assign T1923 = T1382 & T1924;
  assign T1924 = T1770[2'h3:2'h3];
  assign T1925 = T1777 & T1924;
  assign T1926 = {readyToXmit_4_3, readyToXmit_3_3};
  assign readyToXmit_3_3 = T1927;
  assign T1927 = T1931 ? T1790 : T1928;
  assign T1928 = T1929 ? T1782 : 1'h0;
  assign T1929 = T1238 & T1930;
  assign T1930 = T1788[2'h3:2'h3];
  assign T1931 = T1795 & T1930;
  assign readyToXmit_4_3 = T1932;
  assign T1932 = T1936 ? T1807 : T1933;
  assign T1933 = T1934 ? T1799 : 1'h0;
  assign T1934 = T1094 & T1935;
  assign T1935 = T1805[2'h3:2'h3];
  assign T1936 = T1812 & T1935;
  assign T1937 = {T1955, T1938};
  assign T1938 = {readyToXmit_7_3, T1939};
  assign T1939 = {readyToXmit_6_3, readyToXmit_5_3};
  assign readyToXmit_5_3 = T1940;
  assign T1940 = T1944 ? T1827 : T1941;
  assign T1941 = T1942 ? T1819 : 1'h0;
  assign T1942 = T950 & T1943;
  assign T1943 = T1825[2'h3:2'h3];
  assign T1944 = T1832 & T1943;
  assign readyToXmit_6_3 = T1945;
  assign T1945 = T1949 ? T1844 : T1946;
  assign T1946 = T1947 ? T1836 : 1'h0;
  assign T1947 = T806 & T1948;
  assign T1948 = T1842[2'h3:2'h3];
  assign T1949 = T1849 & T1948;
  assign readyToXmit_7_3 = T1950;
  assign T1950 = T1954 ? T1861 : T1951;
  assign T1951 = T1952 ? T1853 : 1'h0;
  assign T1952 = T662 & T1953;
  assign T1953 = T1859[2'h3:2'h3];
  assign T1954 = T1866 & T1953;
  assign T1955 = {readyToXmit_9_3, readyToXmit_8_3};
  assign readyToXmit_8_3 = T1956;
  assign T1956 = T1960 ? T1879 : T1957;
  assign T1957 = T1958 ? T1871 : 1'h0;
  assign T1958 = T518 & T1959;
  assign T1959 = T1877[2'h3:2'h3];
  assign T1960 = T1884 & T1959;
  assign readyToXmit_9_3 = T1961;
  assign T1961 = T1965 ? T1896 : T1962;
  assign T1962 = T1963 ? T1888 : 1'h0;
  assign T1963 = T374 & T1964;
  assign T1964 = T1894[2'h3:2'h3];
  assign T1965 = T1901 & T1964;
  assign T1966 = T1967 ? CreditCon_5_io_outCredit : CreditCon_4_io_outCredit;
  assign T1967 = T246;
  assign T1968 = T1969 != 10'h0;
  assign T1969 = T1970;
  assign T1970 = {T2000, T1971};
  assign T1971 = {T1989, T1972};
  assign T1972 = {readyToXmit_2_2, T1973};
  assign T1973 = {readyToXmit_1_2, readyToXmit_0_2};
  assign readyToXmit_0_2 = T1974;
  assign T1974 = T1978 ? T1738 : T1975;
  assign T1975 = T1976 ? T1730 : 1'h0;
  assign T1976 = T1670 & T1977;
  assign T1977 = T1736[2'h2:2'h2];
  assign T1978 = T1743 & T1977;
  assign readyToXmit_1_2 = T1979;
  assign T1979 = T1983 ? T1755 : T1980;
  assign T1980 = T1981 ? T1747 : 1'h0;
  assign T1981 = T1526 & T1982;
  assign T1982 = T1753[2'h2:2'h2];
  assign T1983 = T1760 & T1982;
  assign readyToXmit_2_2 = T1984;
  assign T1984 = T1988 ? T1772 : T1985;
  assign T1985 = T1986 ? T1764 : 1'h0;
  assign T1986 = T1382 & T1987;
  assign T1987 = T1770[2'h2:2'h2];
  assign T1988 = T1777 & T1987;
  assign T1989 = {readyToXmit_4_2, readyToXmit_3_2};
  assign readyToXmit_3_2 = T1990;
  assign T1990 = T1994 ? T1790 : T1991;
  assign T1991 = T1992 ? T1782 : 1'h0;
  assign T1992 = T1238 & T1993;
  assign T1993 = T1788[2'h2:2'h2];
  assign T1994 = T1795 & T1993;
  assign readyToXmit_4_2 = T1995;
  assign T1995 = T1999 ? T1807 : T1996;
  assign T1996 = T1997 ? T1799 : 1'h0;
  assign T1997 = T1094 & T1998;
  assign T1998 = T1805[2'h2:2'h2];
  assign T1999 = T1812 & T1998;
  assign T2000 = {T2018, T2001};
  assign T2001 = {readyToXmit_7_2, T2002};
  assign T2002 = {readyToXmit_6_2, readyToXmit_5_2};
  assign readyToXmit_5_2 = T2003;
  assign T2003 = T2007 ? T1827 : T2004;
  assign T2004 = T2005 ? T1819 : 1'h0;
  assign T2005 = T950 & T2006;
  assign T2006 = T1825[2'h2:2'h2];
  assign T2007 = T1832 & T2006;
  assign readyToXmit_6_2 = T2008;
  assign T2008 = T2012 ? T1844 : T2009;
  assign T2009 = T2010 ? T1836 : 1'h0;
  assign T2010 = T806 & T2011;
  assign T2011 = T1842[2'h2:2'h2];
  assign T2012 = T1849 & T2011;
  assign readyToXmit_7_2 = T2013;
  assign T2013 = T2017 ? T1861 : T2014;
  assign T2014 = T2015 ? T1853 : 1'h0;
  assign T2015 = T662 & T2016;
  assign T2016 = T1859[2'h2:2'h2];
  assign T2017 = T1866 & T2016;
  assign T2018 = {readyToXmit_9_2, readyToXmit_8_2};
  assign readyToXmit_8_2 = T2019;
  assign T2019 = T2023 ? T1879 : T2020;
  assign T2020 = T2021 ? T1871 : 1'h0;
  assign T2021 = T518 & T2022;
  assign T2022 = T1877[2'h2:2'h2];
  assign T2023 = T1884 & T2022;
  assign readyToXmit_9_2 = T2024;
  assign T2024 = T2028 ? T1896 : T2025;
  assign T2025 = T2026 ? T1888 : 1'h0;
  assign T2026 = T374 & T2027;
  assign T2027 = T1894[2'h2:2'h2];
  assign T2028 = T1901 & T2027;
  assign T2029 = T2030 ? CreditCon_3_io_outCredit : CreditCon_2_io_outCredit;
  assign T2030 = T258;
  assign T2031 = T2032 != 10'h0;
  assign T2032 = T2033;
  assign T2033 = {T2063, T2034};
  assign T2034 = {T2052, T2035};
  assign T2035 = {readyToXmit_2_1, T2036};
  assign T2036 = {readyToXmit_1_1, readyToXmit_0_1};
  assign readyToXmit_0_1 = T2037;
  assign T2037 = T2041 ? T1738 : T2038;
  assign T2038 = T2039 ? T1730 : 1'h0;
  assign T2039 = T1670 & T2040;
  assign T2040 = T1736[1'h1:1'h1];
  assign T2041 = T1743 & T2040;
  assign readyToXmit_1_1 = T2042;
  assign T2042 = T2046 ? T1755 : T2043;
  assign T2043 = T2044 ? T1747 : 1'h0;
  assign T2044 = T1526 & T2045;
  assign T2045 = T1753[1'h1:1'h1];
  assign T2046 = T1760 & T2045;
  assign readyToXmit_2_1 = T2047;
  assign T2047 = T2051 ? T1772 : T2048;
  assign T2048 = T2049 ? T1764 : 1'h0;
  assign T2049 = T1382 & T2050;
  assign T2050 = T1770[1'h1:1'h1];
  assign T2051 = T1777 & T2050;
  assign T2052 = {readyToXmit_4_1, readyToXmit_3_1};
  assign readyToXmit_3_1 = T2053;
  assign T2053 = T2057 ? T1790 : T2054;
  assign T2054 = T2055 ? T1782 : 1'h0;
  assign T2055 = T1238 & T2056;
  assign T2056 = T1788[1'h1:1'h1];
  assign T2057 = T1795 & T2056;
  assign readyToXmit_4_1 = T2058;
  assign T2058 = T2062 ? T1807 : T2059;
  assign T2059 = T2060 ? T1799 : 1'h0;
  assign T2060 = T1094 & T2061;
  assign T2061 = T1805[1'h1:1'h1];
  assign T2062 = T1812 & T2061;
  assign T2063 = {T2081, T2064};
  assign T2064 = {readyToXmit_7_1, T2065};
  assign T2065 = {readyToXmit_6_1, readyToXmit_5_1};
  assign readyToXmit_5_1 = T2066;
  assign T2066 = T2070 ? T1827 : T2067;
  assign T2067 = T2068 ? T1819 : 1'h0;
  assign T2068 = T950 & T2069;
  assign T2069 = T1825[1'h1:1'h1];
  assign T2070 = T1832 & T2069;
  assign readyToXmit_6_1 = T2071;
  assign T2071 = T2075 ? T1844 : T2072;
  assign T2072 = T2073 ? T1836 : 1'h0;
  assign T2073 = T806 & T2074;
  assign T2074 = T1842[1'h1:1'h1];
  assign T2075 = T1849 & T2074;
  assign readyToXmit_7_1 = T2076;
  assign T2076 = T2080 ? T1861 : T2077;
  assign T2077 = T2078 ? T1853 : 1'h0;
  assign T2078 = T662 & T2079;
  assign T2079 = T1859[1'h1:1'h1];
  assign T2080 = T1866 & T2079;
  assign T2081 = {readyToXmit_9_1, readyToXmit_8_1};
  assign readyToXmit_8_1 = T2082;
  assign T2082 = T2086 ? T1879 : T2083;
  assign T2083 = T2084 ? T1871 : 1'h0;
  assign T2084 = T518 & T2085;
  assign T2085 = T1877[1'h1:1'h1];
  assign T2086 = T1884 & T2085;
  assign readyToXmit_9_1 = T2087;
  assign T2087 = T2091 ? T1896 : T2088;
  assign T2088 = T2089 ? T1888 : 1'h0;
  assign T2089 = T374 & T2090;
  assign T2090 = T1894[1'h1:1'h1];
  assign T2091 = T1901 & T2090;
  assign T2092 = T2093 ? CreditCon_1_io_outCredit : CreditCon_io_outCredit;
  assign T2093 = T270;
  assign T2094 = T2095 != 10'h0;
  assign T2095 = T2096;
  assign T2096 = {T2126, T2097};
  assign T2097 = {T2115, T2098};
  assign T2098 = {readyToXmit_2_0, T2099};
  assign T2099 = {readyToXmit_1_0, readyToXmit_0_0};
  assign readyToXmit_0_0 = T2100;
  assign T2100 = T2104 ? T1738 : T2101;
  assign T2101 = T2102 ? T1730 : 1'h0;
  assign T2102 = T1670 & T2103;
  assign T2103 = T1736[1'h0:1'h0];
  assign T2104 = T1743 & T2103;
  assign readyToXmit_1_0 = T2105;
  assign T2105 = T2109 ? T1755 : T2106;
  assign T2106 = T2107 ? T1747 : 1'h0;
  assign T2107 = T1526 & T2108;
  assign T2108 = T1753[1'h0:1'h0];
  assign T2109 = T1760 & T2108;
  assign readyToXmit_2_0 = T2110;
  assign T2110 = T2114 ? T1772 : T2111;
  assign T2111 = T2112 ? T1764 : 1'h0;
  assign T2112 = T1382 & T2113;
  assign T2113 = T1770[1'h0:1'h0];
  assign T2114 = T1777 & T2113;
  assign T2115 = {readyToXmit_4_0, readyToXmit_3_0};
  assign readyToXmit_3_0 = T2116;
  assign T2116 = T2120 ? T1790 : T2117;
  assign T2117 = T2118 ? T1782 : 1'h0;
  assign T2118 = T1238 & T2119;
  assign T2119 = T1788[1'h0:1'h0];
  assign T2120 = T1795 & T2119;
  assign readyToXmit_4_0 = T2121;
  assign T2121 = T2125 ? T1807 : T2122;
  assign T2122 = T2123 ? T1799 : 1'h0;
  assign T2123 = T1094 & T2124;
  assign T2124 = T1805[1'h0:1'h0];
  assign T2125 = T1812 & T2124;
  assign T2126 = {T2144, T2127};
  assign T2127 = {readyToXmit_7_0, T2128};
  assign T2128 = {readyToXmit_6_0, readyToXmit_5_0};
  assign readyToXmit_5_0 = T2129;
  assign T2129 = T2133 ? T1827 : T2130;
  assign T2130 = T2131 ? T1819 : 1'h0;
  assign T2131 = T950 & T2132;
  assign T2132 = T1825[1'h0:1'h0];
  assign T2133 = T1832 & T2132;
  assign readyToXmit_6_0 = T2134;
  assign T2134 = T2138 ? T1844 : T2135;
  assign T2135 = T2136 ? T1836 : 1'h0;
  assign T2136 = T806 & T2137;
  assign T2137 = T1842[1'h0:1'h0];
  assign T2138 = T1849 & T2137;
  assign readyToXmit_7_0 = T2139;
  assign T2139 = T2143 ? T1861 : T2140;
  assign T2140 = T2141 ? T1853 : 1'h0;
  assign T2141 = T662 & T2142;
  assign T2142 = T1859[1'h0:1'h0];
  assign T2143 = T1866 & T2142;
  assign T2144 = {readyToXmit_9_0, readyToXmit_8_0};
  assign readyToXmit_8_0 = T2145;
  assign T2145 = T2149 ? T1879 : T2146;
  assign T2146 = T2147 ? T1871 : 1'h0;
  assign T2147 = T518 & T2148;
  assign T2148 = T1877[1'h0:1'h0];
  assign T2149 = T1884 & T2148;
  assign readyToXmit_9_0 = T2150;
  assign T2150 = T2154 ? T1896 : T2151;
  assign T2151 = T2152 ? T1888 : 1'h0;
  assign T2152 = T374 & T2153;
  assign T2153 = T1894[1'h0:1'h0];
  assign T2154 = T1901 & T2153;
  assign T2155 = RouterBuffer_io_deq_valid & T2156;
  assign T2156 = 3'h2 <= VCRouterStateManagement_io_currentState;
  assign T2157 = RouterBuffer_1_io_deq_valid & T2158;
  assign T2158 = 3'h2 <= VCRouterStateManagement_1_io_currentState;
  assign T2159 = RouterBuffer_2_io_deq_valid & T2160;
  assign T2160 = 3'h2 <= VCRouterStateManagement_2_io_currentState;
  assign T2161 = RouterBuffer_3_io_deq_valid & T2162;
  assign T2162 = 3'h2 <= VCRouterStateManagement_3_io_currentState;
  assign T2163 = RouterBuffer_4_io_deq_valid & T2164;
  assign T2164 = 3'h2 <= VCRouterStateManagement_4_io_currentState;
  assign T2165 = RouterBuffer_5_io_deq_valid & T2166;
  assign T2166 = 3'h2 <= VCRouterStateManagement_5_io_currentState;
  assign T2167 = RouterBuffer_6_io_deq_valid & T2168;
  assign T2168 = 3'h2 <= VCRouterStateManagement_6_io_currentState;
  assign T2169 = RouterBuffer_7_io_deq_valid & T2170;
  assign T2170 = 3'h2 <= VCRouterStateManagement_7_io_currentState;
  assign T2171 = RouterBuffer_8_io_deq_valid & T2172;
  assign T2172 = 3'h2 <= VCRouterStateManagement_8_io_currentState;
  assign T2173 = RouterBuffer_9_io_deq_valid & T2174;
  assign T2174 = 3'h2 <= VCRouterStateManagement_9_io_currentState;
  assign T2175 = validVCs_0_0[1'h0:1'h0];
  assign T2177 = T2179 & T2178;
  assign T2178 = VCRouterOutputStateManagement_io_currentState == 2'h2;
  assign T2179 = flitsAreTail_0 & CreditCon_io_outCredit;
  assign T2180 = validVCs_0_0[1'h1:1'h1];
  assign T2182 = T2184 & T2183;
  assign T2183 = VCRouterOutputStateManagement_io_currentState == 2'h2;
  assign T2184 = flitsAreTail_0 & CreditCon_1_io_outCredit;
  assign T2185 = validVCs_0_1[1'h0:1'h0];
  assign T2187 = T2189 & T2188;
  assign T2188 = VCRouterOutputStateManagement_1_io_currentState == 2'h2;
  assign T2189 = flitsAreTail_0 & CreditCon_2_io_outCredit;
  assign T2190 = validVCs_0_1[1'h1:1'h1];
  assign T2192 = T2194 & T2193;
  assign T2193 = VCRouterOutputStateManagement_1_io_currentState == 2'h2;
  assign T2194 = flitsAreTail_0 & CreditCon_3_io_outCredit;
  assign T2195 = validVCs_0_2[1'h0:1'h0];
  assign T2197 = T2199 & T2198;
  assign T2198 = VCRouterOutputStateManagement_2_io_currentState == 2'h2;
  assign T2199 = flitsAreTail_0 & CreditCon_4_io_outCredit;
  assign T2200 = validVCs_0_2[1'h1:1'h1];
  assign T2202 = T2204 & T2203;
  assign T2203 = VCRouterOutputStateManagement_2_io_currentState == 2'h2;
  assign T2204 = flitsAreTail_0 & CreditCon_5_io_outCredit;
  assign T2205 = validVCs_0_3[1'h0:1'h0];
  assign T2207 = T2209 & T2208;
  assign T2208 = VCRouterOutputStateManagement_3_io_currentState == 2'h2;
  assign T2209 = flitsAreTail_0 & CreditCon_6_io_outCredit;
  assign T2210 = validVCs_0_3[1'h1:1'h1];
  assign T2212 = T2214 & T2213;
  assign T2213 = VCRouterOutputStateManagement_3_io_currentState == 2'h2;
  assign T2214 = flitsAreTail_0 & CreditCon_7_io_outCredit;
  assign T2215 = validVCs_0_4[1'h0:1'h0];
  assign T2217 = T2219 & T2218;
  assign T2218 = VCRouterOutputStateManagement_4_io_currentState == 2'h2;
  assign T2219 = flitsAreTail_0 & CreditCon_8_io_outCredit;
  assign T2220 = validVCs_0_4[1'h1:1'h1];
  assign T2222 = T2224 & T2223;
  assign T2223 = VCRouterOutputStateManagement_4_io_currentState == 2'h2;
  assign T2224 = flitsAreTail_0 & CreditCon_9_io_outCredit;
  assign T2225 = validVCs_1_0[1'h0:1'h0];
  assign T2227 = T2229 & T2228;
  assign T2228 = VCRouterOutputStateManagement_io_currentState == 2'h2;
  assign T2229 = flitsAreTail_1 & CreditCon_io_outCredit;
  assign T2230 = validVCs_1_0[1'h1:1'h1];
  assign T2232 = T2234 & T2233;
  assign T2233 = VCRouterOutputStateManagement_io_currentState == 2'h2;
  assign T2234 = flitsAreTail_1 & CreditCon_1_io_outCredit;
  assign T2235 = validVCs_1_1[1'h0:1'h0];
  assign T2237 = T2239 & T2238;
  assign T2238 = VCRouterOutputStateManagement_1_io_currentState == 2'h2;
  assign T2239 = flitsAreTail_1 & CreditCon_2_io_outCredit;
  assign T2240 = validVCs_1_1[1'h1:1'h1];
  assign T2242 = T2244 & T2243;
  assign T2243 = VCRouterOutputStateManagement_1_io_currentState == 2'h2;
  assign T2244 = flitsAreTail_1 & CreditCon_3_io_outCredit;
  assign T2245 = validVCs_1_2[1'h0:1'h0];
  assign T2247 = T2249 & T2248;
  assign T2248 = VCRouterOutputStateManagement_2_io_currentState == 2'h2;
  assign T2249 = flitsAreTail_1 & CreditCon_4_io_outCredit;
  assign T2250 = validVCs_1_2[1'h1:1'h1];
  assign T2252 = T2254 & T2253;
  assign T2253 = VCRouterOutputStateManagement_2_io_currentState == 2'h2;
  assign T2254 = flitsAreTail_1 & CreditCon_5_io_outCredit;
  assign T2255 = validVCs_1_3[1'h0:1'h0];
  assign T2257 = T2259 & T2258;
  assign T2258 = VCRouterOutputStateManagement_3_io_currentState == 2'h2;
  assign T2259 = flitsAreTail_1 & CreditCon_6_io_outCredit;
  assign T2260 = validVCs_1_3[1'h1:1'h1];
  assign T2262 = T2264 & T2263;
  assign T2263 = VCRouterOutputStateManagement_3_io_currentState == 2'h2;
  assign T2264 = flitsAreTail_1 & CreditCon_7_io_outCredit;
  assign T2265 = validVCs_1_4[1'h0:1'h0];
  assign T2267 = T2269 & T2268;
  assign T2268 = VCRouterOutputStateManagement_4_io_currentState == 2'h2;
  assign T2269 = flitsAreTail_1 & CreditCon_8_io_outCredit;
  assign T2270 = validVCs_1_4[1'h1:1'h1];
  assign T2272 = T2274 & T2273;
  assign T2273 = VCRouterOutputStateManagement_4_io_currentState == 2'h2;
  assign T2274 = flitsAreTail_1 & CreditCon_9_io_outCredit;
  assign T2275 = validVCs_2_0[1'h0:1'h0];
  assign T2277 = T2279 & T2278;
  assign T2278 = VCRouterOutputStateManagement_io_currentState == 2'h2;
  assign T2279 = flitsAreTail_2 & CreditCon_io_outCredit;
  assign T2280 = validVCs_2_0[1'h1:1'h1];
  assign T2282 = T2284 & T2283;
  assign T2283 = VCRouterOutputStateManagement_io_currentState == 2'h2;
  assign T2284 = flitsAreTail_2 & CreditCon_1_io_outCredit;
  assign T2285 = validVCs_2_1[1'h0:1'h0];
  assign T2287 = T2289 & T2288;
  assign T2288 = VCRouterOutputStateManagement_1_io_currentState == 2'h2;
  assign T2289 = flitsAreTail_2 & CreditCon_2_io_outCredit;
  assign T2290 = validVCs_2_1[1'h1:1'h1];
  assign T2292 = T2294 & T2293;
  assign T2293 = VCRouterOutputStateManagement_1_io_currentState == 2'h2;
  assign T2294 = flitsAreTail_2 & CreditCon_3_io_outCredit;
  assign T2295 = validVCs_2_2[1'h0:1'h0];
  assign T2297 = T2299 & T2298;
  assign T2298 = VCRouterOutputStateManagement_2_io_currentState == 2'h2;
  assign T2299 = flitsAreTail_2 & CreditCon_4_io_outCredit;
  assign T2300 = validVCs_2_2[1'h1:1'h1];
  assign T2302 = T2304 & T2303;
  assign T2303 = VCRouterOutputStateManagement_2_io_currentState == 2'h2;
  assign T2304 = flitsAreTail_2 & CreditCon_5_io_outCredit;
  assign T2305 = validVCs_2_3[1'h0:1'h0];
  assign T2307 = T2309 & T2308;
  assign T2308 = VCRouterOutputStateManagement_3_io_currentState == 2'h2;
  assign T2309 = flitsAreTail_2 & CreditCon_6_io_outCredit;
  assign T2310 = validVCs_2_3[1'h1:1'h1];
  assign T2312 = T2314 & T2313;
  assign T2313 = VCRouterOutputStateManagement_3_io_currentState == 2'h2;
  assign T2314 = flitsAreTail_2 & CreditCon_7_io_outCredit;
  assign T2315 = validVCs_2_4[1'h0:1'h0];
  assign T2317 = T2319 & T2318;
  assign T2318 = VCRouterOutputStateManagement_4_io_currentState == 2'h2;
  assign T2319 = flitsAreTail_2 & CreditCon_8_io_outCredit;
  assign T2320 = validVCs_2_4[1'h1:1'h1];
  assign T2322 = T2324 & T2323;
  assign T2323 = VCRouterOutputStateManagement_4_io_currentState == 2'h2;
  assign T2324 = flitsAreTail_2 & CreditCon_9_io_outCredit;
  assign T2325 = validVCs_3_0[1'h0:1'h0];
  assign T2327 = T2329 & T2328;
  assign T2328 = VCRouterOutputStateManagement_io_currentState == 2'h2;
  assign T2329 = flitsAreTail_3 & CreditCon_io_outCredit;
  assign T2330 = validVCs_3_0[1'h1:1'h1];
  assign T2332 = T2334 & T2333;
  assign T2333 = VCRouterOutputStateManagement_io_currentState == 2'h2;
  assign T2334 = flitsAreTail_3 & CreditCon_1_io_outCredit;
  assign T2335 = validVCs_3_1[1'h0:1'h0];
  assign T2337 = T2339 & T2338;
  assign T2338 = VCRouterOutputStateManagement_1_io_currentState == 2'h2;
  assign T2339 = flitsAreTail_3 & CreditCon_2_io_outCredit;
  assign T2340 = validVCs_3_1[1'h1:1'h1];
  assign T2342 = T2344 & T2343;
  assign T2343 = VCRouterOutputStateManagement_1_io_currentState == 2'h2;
  assign T2344 = flitsAreTail_3 & CreditCon_3_io_outCredit;
  assign T2345 = validVCs_3_2[1'h0:1'h0];
  assign T2347 = T2349 & T2348;
  assign T2348 = VCRouterOutputStateManagement_2_io_currentState == 2'h2;
  assign T2349 = flitsAreTail_3 & CreditCon_4_io_outCredit;
  assign T2350 = validVCs_3_2[1'h1:1'h1];
  assign T2352 = T2354 & T2353;
  assign T2353 = VCRouterOutputStateManagement_2_io_currentState == 2'h2;
  assign T2354 = flitsAreTail_3 & CreditCon_5_io_outCredit;
  assign T2355 = validVCs_3_3[1'h0:1'h0];
  assign T2357 = T2359 & T2358;
  assign T2358 = VCRouterOutputStateManagement_3_io_currentState == 2'h2;
  assign T2359 = flitsAreTail_3 & CreditCon_6_io_outCredit;
  assign T2360 = validVCs_3_3[1'h1:1'h1];
  assign T2362 = T2364 & T2363;
  assign T2363 = VCRouterOutputStateManagement_3_io_currentState == 2'h2;
  assign T2364 = flitsAreTail_3 & CreditCon_7_io_outCredit;
  assign T2365 = validVCs_3_4[1'h0:1'h0];
  assign T2367 = T2369 & T2368;
  assign T2368 = VCRouterOutputStateManagement_4_io_currentState == 2'h2;
  assign T2369 = flitsAreTail_3 & CreditCon_8_io_outCredit;
  assign T2370 = validVCs_3_4[1'h1:1'h1];
  assign T2372 = T2374 & T2373;
  assign T2373 = VCRouterOutputStateManagement_4_io_currentState == 2'h2;
  assign T2374 = flitsAreTail_3 & CreditCon_9_io_outCredit;
  assign T2375 = validVCs_4_0[1'h0:1'h0];
  assign T2377 = T2379 & T2378;
  assign T2378 = VCRouterOutputStateManagement_io_currentState == 2'h2;
  assign T2379 = flitsAreTail_4 & CreditCon_io_outCredit;
  assign T2380 = validVCs_4_0[1'h1:1'h1];
  assign T2382 = T2384 & T2383;
  assign T2383 = VCRouterOutputStateManagement_io_currentState == 2'h2;
  assign T2384 = flitsAreTail_4 & CreditCon_1_io_outCredit;
  assign T2385 = validVCs_4_1[1'h0:1'h0];
  assign T2387 = T2389 & T2388;
  assign T2388 = VCRouterOutputStateManagement_1_io_currentState == 2'h2;
  assign T2389 = flitsAreTail_4 & CreditCon_2_io_outCredit;
  assign T2390 = validVCs_4_1[1'h1:1'h1];
  assign T2392 = T2394 & T2393;
  assign T2393 = VCRouterOutputStateManagement_1_io_currentState == 2'h2;
  assign T2394 = flitsAreTail_4 & CreditCon_3_io_outCredit;
  assign T2395 = validVCs_4_2[1'h0:1'h0];
  assign T2397 = T2399 & T2398;
  assign T2398 = VCRouterOutputStateManagement_2_io_currentState == 2'h2;
  assign T2399 = flitsAreTail_4 & CreditCon_4_io_outCredit;
  assign T2400 = validVCs_4_2[1'h1:1'h1];
  assign T2402 = T2404 & T2403;
  assign T2403 = VCRouterOutputStateManagement_2_io_currentState == 2'h2;
  assign T2404 = flitsAreTail_4 & CreditCon_5_io_outCredit;
  assign T2405 = validVCs_4_3[1'h0:1'h0];
  assign T2407 = T2409 & T2408;
  assign T2408 = VCRouterOutputStateManagement_3_io_currentState == 2'h2;
  assign T2409 = flitsAreTail_4 & CreditCon_6_io_outCredit;
  assign T2410 = validVCs_4_3[1'h1:1'h1];
  assign T2412 = T2414 & T2413;
  assign T2413 = VCRouterOutputStateManagement_3_io_currentState == 2'h2;
  assign T2414 = flitsAreTail_4 & CreditCon_7_io_outCredit;
  assign T2415 = validVCs_4_4[1'h0:1'h0];
  assign T2417 = T2419 & T2418;
  assign T2418 = VCRouterOutputStateManagement_4_io_currentState == 2'h2;
  assign T2419 = flitsAreTail_4 & CreditCon_8_io_outCredit;
  assign T2420 = validVCs_4_4[1'h1:1'h1];
  assign T2422 = T2424 & T2423;
  assign T2423 = VCRouterOutputStateManagement_4_io_currentState == 2'h2;
  assign T2424 = flitsAreTail_4 & CreditCon_9_io_outCredit;
  assign T2425 = validVCs_5_0[1'h0:1'h0];
  assign T2427 = T2429 & T2428;
  assign T2428 = VCRouterOutputStateManagement_io_currentState == 2'h2;
  assign T2429 = flitsAreTail_5 & CreditCon_io_outCredit;
  assign T2430 = validVCs_5_0[1'h1:1'h1];
  assign T2432 = T2434 & T2433;
  assign T2433 = VCRouterOutputStateManagement_io_currentState == 2'h2;
  assign T2434 = flitsAreTail_5 & CreditCon_1_io_outCredit;
  assign T2435 = validVCs_5_1[1'h0:1'h0];
  assign T2437 = T2439 & T2438;
  assign T2438 = VCRouterOutputStateManagement_1_io_currentState == 2'h2;
  assign T2439 = flitsAreTail_5 & CreditCon_2_io_outCredit;
  assign T2440 = validVCs_5_1[1'h1:1'h1];
  assign T2442 = T2444 & T2443;
  assign T2443 = VCRouterOutputStateManagement_1_io_currentState == 2'h2;
  assign T2444 = flitsAreTail_5 & CreditCon_3_io_outCredit;
  assign T2445 = validVCs_5_2[1'h0:1'h0];
  assign T2447 = T2449 & T2448;
  assign T2448 = VCRouterOutputStateManagement_2_io_currentState == 2'h2;
  assign T2449 = flitsAreTail_5 & CreditCon_4_io_outCredit;
  assign T2450 = validVCs_5_2[1'h1:1'h1];
  assign T2452 = T2454 & T2453;
  assign T2453 = VCRouterOutputStateManagement_2_io_currentState == 2'h2;
  assign T2454 = flitsAreTail_5 & CreditCon_5_io_outCredit;
  assign T2455 = validVCs_5_3[1'h0:1'h0];
  assign T2457 = T2459 & T2458;
  assign T2458 = VCRouterOutputStateManagement_3_io_currentState == 2'h2;
  assign T2459 = flitsAreTail_5 & CreditCon_6_io_outCredit;
  assign T2460 = validVCs_5_3[1'h1:1'h1];
  assign T2462 = T2464 & T2463;
  assign T2463 = VCRouterOutputStateManagement_3_io_currentState == 2'h2;
  assign T2464 = flitsAreTail_5 & CreditCon_7_io_outCredit;
  assign T2465 = validVCs_5_4[1'h0:1'h0];
  assign T2467 = T2469 & T2468;
  assign T2468 = VCRouterOutputStateManagement_4_io_currentState == 2'h2;
  assign T2469 = flitsAreTail_5 & CreditCon_8_io_outCredit;
  assign T2470 = validVCs_5_4[1'h1:1'h1];
  assign T2472 = T2474 & T2473;
  assign T2473 = VCRouterOutputStateManagement_4_io_currentState == 2'h2;
  assign T2474 = flitsAreTail_5 & CreditCon_9_io_outCredit;
  assign T2475 = validVCs_6_0[1'h0:1'h0];
  assign T2477 = T2479 & T2478;
  assign T2478 = VCRouterOutputStateManagement_io_currentState == 2'h2;
  assign T2479 = flitsAreTail_6 & CreditCon_io_outCredit;
  assign T2480 = validVCs_6_0[1'h1:1'h1];
  assign T2482 = T2484 & T2483;
  assign T2483 = VCRouterOutputStateManagement_io_currentState == 2'h2;
  assign T2484 = flitsAreTail_6 & CreditCon_1_io_outCredit;
  assign T2485 = validVCs_6_1[1'h0:1'h0];
  assign T2487 = T2489 & T2488;
  assign T2488 = VCRouterOutputStateManagement_1_io_currentState == 2'h2;
  assign T2489 = flitsAreTail_6 & CreditCon_2_io_outCredit;
  assign T2490 = validVCs_6_1[1'h1:1'h1];
  assign T2492 = T2494 & T2493;
  assign T2493 = VCRouterOutputStateManagement_1_io_currentState == 2'h2;
  assign T2494 = flitsAreTail_6 & CreditCon_3_io_outCredit;
  assign T2495 = validVCs_6_2[1'h0:1'h0];
  assign T2497 = T2499 & T2498;
  assign T2498 = VCRouterOutputStateManagement_2_io_currentState == 2'h2;
  assign T2499 = flitsAreTail_6 & CreditCon_4_io_outCredit;
  assign T2500 = validVCs_6_2[1'h1:1'h1];
  assign T2502 = T2504 & T2503;
  assign T2503 = VCRouterOutputStateManagement_2_io_currentState == 2'h2;
  assign T2504 = flitsAreTail_6 & CreditCon_5_io_outCredit;
  assign T2505 = validVCs_6_3[1'h0:1'h0];
  assign T2507 = T2509 & T2508;
  assign T2508 = VCRouterOutputStateManagement_3_io_currentState == 2'h2;
  assign T2509 = flitsAreTail_6 & CreditCon_6_io_outCredit;
  assign T2510 = validVCs_6_3[1'h1:1'h1];
  assign T2512 = T2514 & T2513;
  assign T2513 = VCRouterOutputStateManagement_3_io_currentState == 2'h2;
  assign T2514 = flitsAreTail_6 & CreditCon_7_io_outCredit;
  assign T2515 = validVCs_6_4[1'h0:1'h0];
  assign T2517 = T2519 & T2518;
  assign T2518 = VCRouterOutputStateManagement_4_io_currentState == 2'h2;
  assign T2519 = flitsAreTail_6 & CreditCon_8_io_outCredit;
  assign T2520 = validVCs_6_4[1'h1:1'h1];
  assign T2522 = T2524 & T2523;
  assign T2523 = VCRouterOutputStateManagement_4_io_currentState == 2'h2;
  assign T2524 = flitsAreTail_6 & CreditCon_9_io_outCredit;
  assign T2525 = validVCs_7_0[1'h0:1'h0];
  assign T2527 = T2529 & T2528;
  assign T2528 = VCRouterOutputStateManagement_io_currentState == 2'h2;
  assign T2529 = flitsAreTail_7 & CreditCon_io_outCredit;
  assign T2530 = validVCs_7_0[1'h1:1'h1];
  assign T2532 = T2534 & T2533;
  assign T2533 = VCRouterOutputStateManagement_io_currentState == 2'h2;
  assign T2534 = flitsAreTail_7 & CreditCon_1_io_outCredit;
  assign T2535 = validVCs_7_1[1'h0:1'h0];
  assign T2537 = T2539 & T2538;
  assign T2538 = VCRouterOutputStateManagement_1_io_currentState == 2'h2;
  assign T2539 = flitsAreTail_7 & CreditCon_2_io_outCredit;
  assign T2540 = validVCs_7_1[1'h1:1'h1];
  assign T2542 = T2544 & T2543;
  assign T2543 = VCRouterOutputStateManagement_1_io_currentState == 2'h2;
  assign T2544 = flitsAreTail_7 & CreditCon_3_io_outCredit;
  assign T2545 = validVCs_7_2[1'h0:1'h0];
  assign T2547 = T2549 & T2548;
  assign T2548 = VCRouterOutputStateManagement_2_io_currentState == 2'h2;
  assign T2549 = flitsAreTail_7 & CreditCon_4_io_outCredit;
  assign T2550 = validVCs_7_2[1'h1:1'h1];
  assign T2552 = T2554 & T2553;
  assign T2553 = VCRouterOutputStateManagement_2_io_currentState == 2'h2;
  assign T2554 = flitsAreTail_7 & CreditCon_5_io_outCredit;
  assign T2555 = validVCs_7_3[1'h0:1'h0];
  assign T2557 = T2559 & T2558;
  assign T2558 = VCRouterOutputStateManagement_3_io_currentState == 2'h2;
  assign T2559 = flitsAreTail_7 & CreditCon_6_io_outCredit;
  assign T2560 = validVCs_7_3[1'h1:1'h1];
  assign T2562 = T2564 & T2563;
  assign T2563 = VCRouterOutputStateManagement_3_io_currentState == 2'h2;
  assign T2564 = flitsAreTail_7 & CreditCon_7_io_outCredit;
  assign T2565 = validVCs_7_4[1'h0:1'h0];
  assign T2567 = T2569 & T2568;
  assign T2568 = VCRouterOutputStateManagement_4_io_currentState == 2'h2;
  assign T2569 = flitsAreTail_7 & CreditCon_8_io_outCredit;
  assign T2570 = validVCs_7_4[1'h1:1'h1];
  assign T2572 = T2574 & T2573;
  assign T2573 = VCRouterOutputStateManagement_4_io_currentState == 2'h2;
  assign T2574 = flitsAreTail_7 & CreditCon_9_io_outCredit;
  assign T2575 = validVCs_8_0[1'h0:1'h0];
  assign T2577 = T2579 & T2578;
  assign T2578 = VCRouterOutputStateManagement_io_currentState == 2'h2;
  assign T2579 = flitsAreTail_8 & CreditCon_io_outCredit;
  assign T2580 = validVCs_8_0[1'h1:1'h1];
  assign T2582 = T2584 & T2583;
  assign T2583 = VCRouterOutputStateManagement_io_currentState == 2'h2;
  assign T2584 = flitsAreTail_8 & CreditCon_1_io_outCredit;
  assign T2585 = validVCs_8_1[1'h0:1'h0];
  assign T2587 = T2589 & T2588;
  assign T2588 = VCRouterOutputStateManagement_1_io_currentState == 2'h2;
  assign T2589 = flitsAreTail_8 & CreditCon_2_io_outCredit;
  assign T2590 = validVCs_8_1[1'h1:1'h1];
  assign T2592 = T2594 & T2593;
  assign T2593 = VCRouterOutputStateManagement_1_io_currentState == 2'h2;
  assign T2594 = flitsAreTail_8 & CreditCon_3_io_outCredit;
  assign T2595 = validVCs_8_2[1'h0:1'h0];
  assign T2597 = T2599 & T2598;
  assign T2598 = VCRouterOutputStateManagement_2_io_currentState == 2'h2;
  assign T2599 = flitsAreTail_8 & CreditCon_4_io_outCredit;
  assign T2600 = validVCs_8_2[1'h1:1'h1];
  assign T2602 = T2604 & T2603;
  assign T2603 = VCRouterOutputStateManagement_2_io_currentState == 2'h2;
  assign T2604 = flitsAreTail_8 & CreditCon_5_io_outCredit;
  assign T2605 = validVCs_8_3[1'h0:1'h0];
  assign T2607 = T2609 & T2608;
  assign T2608 = VCRouterOutputStateManagement_3_io_currentState == 2'h2;
  assign T2609 = flitsAreTail_8 & CreditCon_6_io_outCredit;
  assign T2610 = validVCs_8_3[1'h1:1'h1];
  assign T2612 = T2614 & T2613;
  assign T2613 = VCRouterOutputStateManagement_3_io_currentState == 2'h2;
  assign T2614 = flitsAreTail_8 & CreditCon_7_io_outCredit;
  assign T2615 = validVCs_8_4[1'h0:1'h0];
  assign T2617 = T2619 & T2618;
  assign T2618 = VCRouterOutputStateManagement_4_io_currentState == 2'h2;
  assign T2619 = flitsAreTail_8 & CreditCon_8_io_outCredit;
  assign T2620 = validVCs_8_4[1'h1:1'h1];
  assign T2622 = T2624 & T2623;
  assign T2623 = VCRouterOutputStateManagement_4_io_currentState == 2'h2;
  assign T2624 = flitsAreTail_8 & CreditCon_9_io_outCredit;
  assign T2625 = validVCs_9_0[1'h0:1'h0];
  assign T2627 = T2629 & T2628;
  assign T2628 = VCRouterOutputStateManagement_io_currentState == 2'h2;
  assign T2629 = flitsAreTail_9 & CreditCon_io_outCredit;
  assign T2630 = validVCs_9_0[1'h1:1'h1];
  assign T2632 = T2634 & T2633;
  assign T2633 = VCRouterOutputStateManagement_io_currentState == 2'h2;
  assign T2634 = flitsAreTail_9 & CreditCon_1_io_outCredit;
  assign T2635 = validVCs_9_1[1'h0:1'h0];
  assign T2637 = T2639 & T2638;
  assign T2638 = VCRouterOutputStateManagement_1_io_currentState == 2'h2;
  assign T2639 = flitsAreTail_9 & CreditCon_2_io_outCredit;
  assign T2640 = validVCs_9_1[1'h1:1'h1];
  assign T2642 = T2644 & T2643;
  assign T2643 = VCRouterOutputStateManagement_1_io_currentState == 2'h2;
  assign T2644 = flitsAreTail_9 & CreditCon_3_io_outCredit;
  assign T2645 = validVCs_9_2[1'h0:1'h0];
  assign T2647 = T2649 & T2648;
  assign T2648 = VCRouterOutputStateManagement_2_io_currentState == 2'h2;
  assign T2649 = flitsAreTail_9 & CreditCon_4_io_outCredit;
  assign T2650 = validVCs_9_2[1'h1:1'h1];
  assign T2652 = T2654 & T2653;
  assign T2653 = VCRouterOutputStateManagement_2_io_currentState == 2'h2;
  assign T2654 = flitsAreTail_9 & CreditCon_5_io_outCredit;
  assign T2655 = validVCs_9_3[1'h0:1'h0];
  assign T2657 = T2659 & T2658;
  assign T2658 = VCRouterOutputStateManagement_3_io_currentState == 2'h2;
  assign T2659 = flitsAreTail_9 & CreditCon_6_io_outCredit;
  assign T2660 = validVCs_9_3[1'h1:1'h1];
  assign T2662 = T2664 & T2663;
  assign T2663 = VCRouterOutputStateManagement_3_io_currentState == 2'h2;
  assign T2664 = flitsAreTail_9 & CreditCon_7_io_outCredit;
  assign T2665 = validVCs_9_4[1'h0:1'h0];
  assign T2667 = T2669 & T2668;
  assign T2668 = VCRouterOutputStateManagement_4_io_currentState == 2'h2;
  assign T2669 = flitsAreTail_9 & CreditCon_8_io_outCredit;
  assign T2670 = validVCs_9_4[1'h1:1'h1];
  assign T2672 = T2674 & T2673;
  assign T2673 = VCRouterOutputStateManagement_4_io_currentState == 2'h2;
  assign T2674 = flitsAreTail_9 & CreditCon_9_io_outCredit;
  assign T3182 = reset ? 3'h0 : T2676;
  assign T2676 = T1670 ? T2677 : R2675;
  assign T2677 = T2678[2'h2:1'h0];
  assign T2678 = RouterBuffer_io_deq_bits_x[5'h1f:1'h1];
  assign T2679 = T2681 & T2680;
  assign T2680 = 3'h3 <= VCRouterStateManagement_io_currentState;
  assign T2681 = T2682;
  assign T2682 = R2683[1'h0:1'h0];
  assign T3183 = reset ? 8'h0 : T2684;
  assign T2684 = 1'h1 << CMeshDOR_io_result;
  assign T2685 = T2687 & T2686;
  assign T2686 = VCRouterStateManagement_io_currentState == 3'h4;
  assign T2687 = R2688;
  assign T3184 = reset ? 1'h1 : T1692;
  assign T3185 = reset ? 3'h0 : T2690;
  assign T2690 = T1526 ? T2691 : R2689;
  assign T2691 = T2692[2'h2:1'h0];
  assign T2692 = RouterBuffer_1_io_deq_bits_x[5'h1f:1'h1];
  assign T2693 = T2695 & T2694;
  assign T2694 = 3'h3 <= VCRouterStateManagement_1_io_currentState;
  assign T2695 = T2696;
  assign T2696 = R2697[1'h0:1'h0];
  assign T3186 = reset ? 8'h0 : T2698;
  assign T2698 = 1'h1 << CMeshDOR_1_io_result;
  assign T2699 = T2701 & T2700;
  assign T2700 = VCRouterStateManagement_1_io_currentState == 3'h4;
  assign T2701 = R2702;
  assign T3187 = reset ? 1'h1 : T1548;
  assign T3188 = reset ? 3'h0 : T2704;
  assign T2704 = T1382 ? T2705 : R2703;
  assign T2705 = T2706[2'h2:1'h0];
  assign T2706 = RouterBuffer_2_io_deq_bits_x[5'h1f:1'h1];
  assign T2707 = T2709 & T2708;
  assign T2708 = 3'h3 <= VCRouterStateManagement_2_io_currentState;
  assign T2709 = T2710;
  assign T2710 = R2711[1'h0:1'h0];
  assign T3189 = reset ? 8'h0 : T2712;
  assign T2712 = 1'h1 << CMeshDOR_2_io_result;
  assign T2713 = T2715 & T2714;
  assign T2714 = VCRouterStateManagement_2_io_currentState == 3'h4;
  assign T2715 = R2716;
  assign T3190 = reset ? 1'h1 : T1404;
  assign T3191 = reset ? 3'h0 : T2718;
  assign T2718 = T1238 ? T2719 : R2717;
  assign T2719 = T2720[2'h2:1'h0];
  assign T2720 = RouterBuffer_3_io_deq_bits_x[5'h1f:1'h1];
  assign T2721 = T2723 & T2722;
  assign T2722 = 3'h3 <= VCRouterStateManagement_3_io_currentState;
  assign T2723 = T2724;
  assign T2724 = R2725[1'h0:1'h0];
  assign T3192 = reset ? 8'h0 : T2726;
  assign T2726 = 1'h1 << CMeshDOR_3_io_result;
  assign T2727 = T2729 & T2728;
  assign T2728 = VCRouterStateManagement_3_io_currentState == 3'h4;
  assign T2729 = R2730;
  assign T3193 = reset ? 1'h1 : T1260;
  assign T3194 = reset ? 3'h0 : T2732;
  assign T2732 = T1094 ? T2733 : R2731;
  assign T2733 = T2734[2'h2:1'h0];
  assign T2734 = RouterBuffer_4_io_deq_bits_x[5'h1f:1'h1];
  assign T2735 = T2737 & T2736;
  assign T2736 = 3'h3 <= VCRouterStateManagement_4_io_currentState;
  assign T2737 = T2738;
  assign T2738 = R2739[1'h0:1'h0];
  assign T3195 = reset ? 8'h0 : T2740;
  assign T2740 = 1'h1 << CMeshDOR_4_io_result;
  assign T2741 = T2743 & T2742;
  assign T2742 = VCRouterStateManagement_4_io_currentState == 3'h4;
  assign T2743 = R2744;
  assign T3196 = reset ? 1'h1 : T1116;
  assign T3197 = reset ? 3'h0 : T2746;
  assign T2746 = T950 ? T2747 : R2745;
  assign T2747 = T2748[2'h2:1'h0];
  assign T2748 = RouterBuffer_5_io_deq_bits_x[5'h1f:1'h1];
  assign T2749 = T2751 & T2750;
  assign T2750 = 3'h3 <= VCRouterStateManagement_5_io_currentState;
  assign T2751 = T2752;
  assign T2752 = R2753[1'h0:1'h0];
  assign T3198 = reset ? 8'h0 : T2754;
  assign T2754 = 1'h1 << CMeshDOR_5_io_result;
  assign T2755 = T2757 & T2756;
  assign T2756 = VCRouterStateManagement_5_io_currentState == 3'h4;
  assign T2757 = R2758;
  assign T3199 = reset ? 1'h1 : T972;
  assign T3200 = reset ? 3'h0 : T2760;
  assign T2760 = T806 ? T2761 : R2759;
  assign T2761 = T2762[2'h2:1'h0];
  assign T2762 = RouterBuffer_6_io_deq_bits_x[5'h1f:1'h1];
  assign T2763 = T2765 & T2764;
  assign T2764 = 3'h3 <= VCRouterStateManagement_6_io_currentState;
  assign T2765 = T2766;
  assign T2766 = R2767[1'h0:1'h0];
  assign T3201 = reset ? 8'h0 : T2768;
  assign T2768 = 1'h1 << CMeshDOR_6_io_result;
  assign T2769 = T2771 & T2770;
  assign T2770 = VCRouterStateManagement_6_io_currentState == 3'h4;
  assign T2771 = R2772;
  assign T3202 = reset ? 1'h1 : T828;
  assign T3203 = reset ? 3'h0 : T2774;
  assign T2774 = T662 ? T2775 : R2773;
  assign T2775 = T2776[2'h2:1'h0];
  assign T2776 = RouterBuffer_7_io_deq_bits_x[5'h1f:1'h1];
  assign T2777 = T2779 & T2778;
  assign T2778 = 3'h3 <= VCRouterStateManagement_7_io_currentState;
  assign T2779 = T2780;
  assign T2780 = R2781[1'h0:1'h0];
  assign T3204 = reset ? 8'h0 : T2782;
  assign T2782 = 1'h1 << CMeshDOR_7_io_result;
  assign T2783 = T2785 & T2784;
  assign T2784 = VCRouterStateManagement_7_io_currentState == 3'h4;
  assign T2785 = R2786;
  assign T3205 = reset ? 1'h1 : T684;
  assign T3206 = reset ? 3'h0 : T2788;
  assign T2788 = T518 ? T2789 : R2787;
  assign T2789 = T2790[2'h2:1'h0];
  assign T2790 = RouterBuffer_8_io_deq_bits_x[5'h1f:1'h1];
  assign T2791 = T2793 & T2792;
  assign T2792 = 3'h3 <= VCRouterStateManagement_8_io_currentState;
  assign T2793 = T2794;
  assign T2794 = R2795[1'h0:1'h0];
  assign T3207 = reset ? 8'h0 : T2796;
  assign T2796 = 1'h1 << CMeshDOR_8_io_result;
  assign T2797 = T2799 & T2798;
  assign T2798 = VCRouterStateManagement_8_io_currentState == 3'h4;
  assign T2799 = R2800;
  assign T3208 = reset ? 1'h1 : T540;
  assign T3209 = reset ? 3'h0 : T2802;
  assign T2802 = T374 ? T2803 : R2801;
  assign T2803 = T2804[2'h2:1'h0];
  assign T2804 = RouterBuffer_9_io_deq_bits_x[5'h1f:1'h1];
  assign T2805 = T2807 & T2806;
  assign T2806 = 3'h3 <= VCRouterStateManagement_9_io_currentState;
  assign T2807 = T2808;
  assign T2808 = R2809[1'h0:1'h0];
  assign T3210 = reset ? 8'h0 : T2810;
  assign T2810 = 1'h1 << CMeshDOR_9_io_result;
  assign T2811 = T2813 & T2812;
  assign T2812 = VCRouterStateManagement_9_io_currentState == 3'h4;
  assign T2813 = R2814;
  assign T3211 = reset ? 1'h1 : T396;
  assign T2815 = T2817 & T2816;
  assign T2816 = 3'h3 <= VCRouterStateManagement_io_currentState;
  assign T2817 = T2818;
  assign T2818 = R2683[1'h1:1'h1];
  assign T2819 = T2821 & T2820;
  assign T2820 = VCRouterStateManagement_io_currentState == 3'h4;
  assign T2821 = R2688;
  assign T2822 = T2824 & T2823;
  assign T2823 = 3'h3 <= VCRouterStateManagement_1_io_currentState;
  assign T2824 = T2825;
  assign T2825 = R2697[1'h1:1'h1];
  assign T2826 = T2828 & T2827;
  assign T2827 = VCRouterStateManagement_1_io_currentState == 3'h4;
  assign T2828 = R2702;
  assign T2829 = T2831 & T2830;
  assign T2830 = 3'h3 <= VCRouterStateManagement_2_io_currentState;
  assign T2831 = T2832;
  assign T2832 = R2711[1'h1:1'h1];
  assign T2833 = T2835 & T2834;
  assign T2834 = VCRouterStateManagement_2_io_currentState == 3'h4;
  assign T2835 = R2716;
  assign T2836 = T2838 & T2837;
  assign T2837 = 3'h3 <= VCRouterStateManagement_3_io_currentState;
  assign T2838 = T2839;
  assign T2839 = R2725[1'h1:1'h1];
  assign T2840 = T2842 & T2841;
  assign T2841 = VCRouterStateManagement_3_io_currentState == 3'h4;
  assign T2842 = R2730;
  assign T2843 = T2845 & T2844;
  assign T2844 = 3'h3 <= VCRouterStateManagement_4_io_currentState;
  assign T2845 = T2846;
  assign T2846 = R2739[1'h1:1'h1];
  assign T2847 = T2849 & T2848;
  assign T2848 = VCRouterStateManagement_4_io_currentState == 3'h4;
  assign T2849 = R2744;
  assign T2850 = T2852 & T2851;
  assign T2851 = 3'h3 <= VCRouterStateManagement_5_io_currentState;
  assign T2852 = T2853;
  assign T2853 = R2753[1'h1:1'h1];
  assign T2854 = T2856 & T2855;
  assign T2855 = VCRouterStateManagement_5_io_currentState == 3'h4;
  assign T2856 = R2758;
  assign T2857 = T2859 & T2858;
  assign T2858 = 3'h3 <= VCRouterStateManagement_6_io_currentState;
  assign T2859 = T2860;
  assign T2860 = R2767[1'h1:1'h1];
  assign T2861 = T2863 & T2862;
  assign T2862 = VCRouterStateManagement_6_io_currentState == 3'h4;
  assign T2863 = R2772;
  assign T2864 = T2866 & T2865;
  assign T2865 = 3'h3 <= VCRouterStateManagement_7_io_currentState;
  assign T2866 = T2867;
  assign T2867 = R2781[1'h1:1'h1];
  assign T2868 = T2870 & T2869;
  assign T2869 = VCRouterStateManagement_7_io_currentState == 3'h4;
  assign T2870 = R2786;
  assign T2871 = T2873 & T2872;
  assign T2872 = 3'h3 <= VCRouterStateManagement_8_io_currentState;
  assign T2873 = T2874;
  assign T2874 = R2795[1'h1:1'h1];
  assign T2875 = T2877 & T2876;
  assign T2876 = VCRouterStateManagement_8_io_currentState == 3'h4;
  assign T2877 = R2800;
  assign T2878 = T2880 & T2879;
  assign T2879 = 3'h3 <= VCRouterStateManagement_9_io_currentState;
  assign T2880 = T2881;
  assign T2881 = R2809[1'h1:1'h1];
  assign T2882 = T2884 & T2883;
  assign T2883 = VCRouterStateManagement_9_io_currentState == 3'h4;
  assign T2884 = R2814;
  assign T2885 = T2887 & T2886;
  assign T2886 = 3'h3 <= VCRouterStateManagement_io_currentState;
  assign T2887 = T2888;
  assign T2888 = R2683[2'h2:2'h2];
  assign T2889 = T2891 & T2890;
  assign T2890 = VCRouterStateManagement_io_currentState == 3'h4;
  assign T2891 = R2688;
  assign T2892 = T2894 & T2893;
  assign T2893 = 3'h3 <= VCRouterStateManagement_1_io_currentState;
  assign T2894 = T2895;
  assign T2895 = R2697[2'h2:2'h2];
  assign T2896 = T2898 & T2897;
  assign T2897 = VCRouterStateManagement_1_io_currentState == 3'h4;
  assign T2898 = R2702;
  assign T2899 = T2901 & T2900;
  assign T2900 = 3'h3 <= VCRouterStateManagement_2_io_currentState;
  assign T2901 = T2902;
  assign T2902 = R2711[2'h2:2'h2];
  assign T2903 = T2905 & T2904;
  assign T2904 = VCRouterStateManagement_2_io_currentState == 3'h4;
  assign T2905 = R2716;
  assign T2906 = T2908 & T2907;
  assign T2907 = 3'h3 <= VCRouterStateManagement_3_io_currentState;
  assign T2908 = T2909;
  assign T2909 = R2725[2'h2:2'h2];
  assign T2910 = T2912 & T2911;
  assign T2911 = VCRouterStateManagement_3_io_currentState == 3'h4;
  assign T2912 = R2730;
  assign T2913 = T2915 & T2914;
  assign T2914 = 3'h3 <= VCRouterStateManagement_4_io_currentState;
  assign T2915 = T2916;
  assign T2916 = R2739[2'h2:2'h2];
  assign T2917 = T2919 & T2918;
  assign T2918 = VCRouterStateManagement_4_io_currentState == 3'h4;
  assign T2919 = R2744;
  assign T2920 = T2922 & T2921;
  assign T2921 = 3'h3 <= VCRouterStateManagement_5_io_currentState;
  assign T2922 = T2923;
  assign T2923 = R2753[2'h2:2'h2];
  assign T2924 = T2926 & T2925;
  assign T2925 = VCRouterStateManagement_5_io_currentState == 3'h4;
  assign T2926 = R2758;
  assign T2927 = T2929 & T2928;
  assign T2928 = 3'h3 <= VCRouterStateManagement_6_io_currentState;
  assign T2929 = T2930;
  assign T2930 = R2767[2'h2:2'h2];
  assign T2931 = T2933 & T2932;
  assign T2932 = VCRouterStateManagement_6_io_currentState == 3'h4;
  assign T2933 = R2772;
  assign T2934 = T2936 & T2935;
  assign T2935 = 3'h3 <= VCRouterStateManagement_7_io_currentState;
  assign T2936 = T2937;
  assign T2937 = R2781[2'h2:2'h2];
  assign T2938 = T2940 & T2939;
  assign T2939 = VCRouterStateManagement_7_io_currentState == 3'h4;
  assign T2940 = R2786;
  assign T2941 = T2943 & T2942;
  assign T2942 = 3'h3 <= VCRouterStateManagement_8_io_currentState;
  assign T2943 = T2944;
  assign T2944 = R2795[2'h2:2'h2];
  assign T2945 = T2947 & T2946;
  assign T2946 = VCRouterStateManagement_8_io_currentState == 3'h4;
  assign T2947 = R2800;
  assign T2948 = T2950 & T2949;
  assign T2949 = 3'h3 <= VCRouterStateManagement_9_io_currentState;
  assign T2950 = T2951;
  assign T2951 = R2809[2'h2:2'h2];
  assign T2952 = T2954 & T2953;
  assign T2953 = VCRouterStateManagement_9_io_currentState == 3'h4;
  assign T2954 = R2814;
  assign T2955 = T2957 & T2956;
  assign T2956 = 3'h3 <= VCRouterStateManagement_io_currentState;
  assign T2957 = T2958;
  assign T2958 = R2683[2'h3:2'h3];
  assign T2959 = T2961 & T2960;
  assign T2960 = VCRouterStateManagement_io_currentState == 3'h4;
  assign T2961 = R2688;
  assign T2962 = T2964 & T2963;
  assign T2963 = 3'h3 <= VCRouterStateManagement_1_io_currentState;
  assign T2964 = T2965;
  assign T2965 = R2697[2'h3:2'h3];
  assign T2966 = T2968 & T2967;
  assign T2967 = VCRouterStateManagement_1_io_currentState == 3'h4;
  assign T2968 = R2702;
  assign T2969 = T2971 & T2970;
  assign T2970 = 3'h3 <= VCRouterStateManagement_2_io_currentState;
  assign T2971 = T2972;
  assign T2972 = R2711[2'h3:2'h3];
  assign T2973 = T2975 & T2974;
  assign T2974 = VCRouterStateManagement_2_io_currentState == 3'h4;
  assign T2975 = R2716;
  assign T2976 = T2978 & T2977;
  assign T2977 = 3'h3 <= VCRouterStateManagement_3_io_currentState;
  assign T2978 = T2979;
  assign T2979 = R2725[2'h3:2'h3];
  assign T2980 = T2982 & T2981;
  assign T2981 = VCRouterStateManagement_3_io_currentState == 3'h4;
  assign T2982 = R2730;
  assign T2983 = T2985 & T2984;
  assign T2984 = 3'h3 <= VCRouterStateManagement_4_io_currentState;
  assign T2985 = T2986;
  assign T2986 = R2739[2'h3:2'h3];
  assign T2987 = T2989 & T2988;
  assign T2988 = VCRouterStateManagement_4_io_currentState == 3'h4;
  assign T2989 = R2744;
  assign T2990 = T2992 & T2991;
  assign T2991 = 3'h3 <= VCRouterStateManagement_5_io_currentState;
  assign T2992 = T2993;
  assign T2993 = R2753[2'h3:2'h3];
  assign T2994 = T2996 & T2995;
  assign T2995 = VCRouterStateManagement_5_io_currentState == 3'h4;
  assign T2996 = R2758;
  assign T2997 = T2999 & T2998;
  assign T2998 = 3'h3 <= VCRouterStateManagement_6_io_currentState;
  assign T2999 = T3000;
  assign T3000 = R2767[2'h3:2'h3];
  assign T3001 = T3003 & T3002;
  assign T3002 = VCRouterStateManagement_6_io_currentState == 3'h4;
  assign T3003 = R2772;
  assign T3004 = T3006 & T3005;
  assign T3005 = 3'h3 <= VCRouterStateManagement_7_io_currentState;
  assign T3006 = T3007;
  assign T3007 = R2781[2'h3:2'h3];
  assign T3008 = T3010 & T3009;
  assign T3009 = VCRouterStateManagement_7_io_currentState == 3'h4;
  assign T3010 = R2786;
  assign T3011 = T3013 & T3012;
  assign T3012 = 3'h3 <= VCRouterStateManagement_8_io_currentState;
  assign T3013 = T3014;
  assign T3014 = R2795[2'h3:2'h3];
  assign T3015 = T3017 & T3016;
  assign T3016 = VCRouterStateManagement_8_io_currentState == 3'h4;
  assign T3017 = R2800;
  assign T3018 = T3020 & T3019;
  assign T3019 = 3'h3 <= VCRouterStateManagement_9_io_currentState;
  assign T3020 = T3021;
  assign T3021 = R2809[2'h3:2'h3];
  assign T3022 = T3024 & T3023;
  assign T3023 = VCRouterStateManagement_9_io_currentState == 3'h4;
  assign T3024 = R2814;
  assign T3025 = T3027 & T3026;
  assign T3026 = 3'h3 <= VCRouterStateManagement_io_currentState;
  assign T3027 = T3028;
  assign T3028 = R2683[3'h4:3'h4];
  assign T3029 = T3031 & T3030;
  assign T3030 = VCRouterStateManagement_io_currentState == 3'h4;
  assign T3031 = R2688;
  assign T3032 = T3034 & T3033;
  assign T3033 = 3'h3 <= VCRouterStateManagement_1_io_currentState;
  assign T3034 = T3035;
  assign T3035 = R2697[3'h4:3'h4];
  assign T3036 = T3038 & T3037;
  assign T3037 = VCRouterStateManagement_1_io_currentState == 3'h4;
  assign T3038 = R2702;
  assign T3039 = T3041 & T3040;
  assign T3040 = 3'h3 <= VCRouterStateManagement_2_io_currentState;
  assign T3041 = T3042;
  assign T3042 = R2711[3'h4:3'h4];
  assign T3043 = T3045 & T3044;
  assign T3044 = VCRouterStateManagement_2_io_currentState == 3'h4;
  assign T3045 = R2716;
  assign T3046 = T3048 & T3047;
  assign T3047 = 3'h3 <= VCRouterStateManagement_3_io_currentState;
  assign T3048 = T3049;
  assign T3049 = R2725[3'h4:3'h4];
  assign T3050 = T3052 & T3051;
  assign T3051 = VCRouterStateManagement_3_io_currentState == 3'h4;
  assign T3052 = R2730;
  assign T3053 = T3055 & T3054;
  assign T3054 = 3'h3 <= VCRouterStateManagement_4_io_currentState;
  assign T3055 = T3056;
  assign T3056 = R2739[3'h4:3'h4];
  assign T3057 = T3059 & T3058;
  assign T3058 = VCRouterStateManagement_4_io_currentState == 3'h4;
  assign T3059 = R2744;
  assign T3060 = T3062 & T3061;
  assign T3061 = 3'h3 <= VCRouterStateManagement_5_io_currentState;
  assign T3062 = T3063;
  assign T3063 = R2753[3'h4:3'h4];
  assign T3064 = T3066 & T3065;
  assign T3065 = VCRouterStateManagement_5_io_currentState == 3'h4;
  assign T3066 = R2758;
  assign T3067 = T3069 & T3068;
  assign T3068 = 3'h3 <= VCRouterStateManagement_6_io_currentState;
  assign T3069 = T3070;
  assign T3070 = R2767[3'h4:3'h4];
  assign T3071 = T3073 & T3072;
  assign T3072 = VCRouterStateManagement_6_io_currentState == 3'h4;
  assign T3073 = R2772;
  assign T3074 = T3076 & T3075;
  assign T3075 = 3'h3 <= VCRouterStateManagement_7_io_currentState;
  assign T3076 = T3077;
  assign T3077 = R2781[3'h4:3'h4];
  assign T3078 = T3080 & T3079;
  assign T3079 = VCRouterStateManagement_7_io_currentState == 3'h4;
  assign T3080 = R2786;
  assign T3081 = T3083 & T3082;
  assign T3082 = 3'h3 <= VCRouterStateManagement_8_io_currentState;
  assign T3083 = T3084;
  assign T3084 = R2795[3'h4:3'h4];
  assign T3085 = T3087 & T3086;
  assign T3086 = VCRouterStateManagement_8_io_currentState == 3'h4;
  assign T3087 = R2800;
  assign T3088 = T3090 & T3089;
  assign T3089 = 3'h3 <= VCRouterStateManagement_9_io_currentState;
  assign T3090 = T3091;
  assign T3091 = R2809[3'h4:3'h4];
  assign T3092 = T3094 & T3093;
  assign T3093 = VCRouterStateManagement_9_io_currentState == 3'h4;
  assign T3094 = R2814;
  assign io_counters_0_counterVal = T3212;
  assign T3212 = {31'h0, T3095};
  assign T3095 = T3096 == 1'h0;
  assign T3096 = T365 ^ 1'h1;
  assign io_outChannels_0_flitValid = R3097;
  assign io_outChannels_0_flit_x = R3098;
  assign T3099 = 55'h0;
  assign T3213 = reset ? T3099 : switch_io_outPorts_0_x;
  assign io_outChannels_1_flitValid = R3100;
  assign io_outChannels_1_flit_x = R3101;
  assign T3102 = 55'h0;
  assign T3214 = reset ? T3102 : switch_io_outPorts_1_x;
  assign io_outChannels_2_flitValid = R3103;
  assign io_outChannels_2_flit_x = R3104;
  assign T3105 = 55'h0;
  assign T3215 = reset ? T3105 : switch_io_outPorts_2_x;
  assign io_outChannels_3_flitValid = R3106;
  assign io_outChannels_3_flit_x = R3107;
  assign T3108 = 55'h0;
  assign T3216 = reset ? T3108 : switch_io_outPorts_3_x;
  assign io_outChannels_4_flitValid = R3109;
  assign io_outChannels_4_flit_x = R3110;
  assign T3111 = 55'h0;
  assign T3217 = reset ? T3111 : switch_io_outPorts_4_x;
  assign io_inChannels_0_credit_0_grant = CreditGen_io_outCredit_grant;
  assign io_inChannels_0_credit_1_grant = CreditGen_1_io_outCredit_grant;
  assign io_inChannels_1_credit_0_grant = CreditGen_2_io_outCredit_grant;
  assign io_inChannels_1_credit_1_grant = CreditGen_3_io_outCredit_grant;
  assign io_inChannels_2_credit_0_grant = CreditGen_4_io_outCredit_grant;
  assign io_inChannels_2_credit_1_grant = CreditGen_5_io_outCredit_grant;
  assign io_inChannels_3_credit_0_grant = CreditGen_6_io_outCredit_grant;
  assign io_inChannels_3_credit_1_grant = CreditGen_7_io_outCredit_grant;
  assign io_inChannels_4_credit_0_grant = CreditGen_8_io_outCredit_grant;
  assign io_inChannels_4_credit_1_grant = CreditGen_9_io_outCredit_grant;
  Switch switch(
       .io_inPorts_9_x( ReplaceVCPort_9_io_newFlit_x ),
       .io_inPorts_8_x( ReplaceVCPort_8_io_newFlit_x ),
       .io_inPorts_7_x( ReplaceVCPort_7_io_newFlit_x ),
       .io_inPorts_6_x( ReplaceVCPort_6_io_newFlit_x ),
       .io_inPorts_5_x( ReplaceVCPort_5_io_newFlit_x ),
       .io_inPorts_4_x( ReplaceVCPort_4_io_newFlit_x ),
       .io_inPorts_3_x( ReplaceVCPort_3_io_newFlit_x ),
       .io_inPorts_2_x( ReplaceVCPort_2_io_newFlit_x ),
       .io_inPorts_1_x( ReplaceVCPort_1_io_newFlit_x ),
       .io_inPorts_0_x( ReplaceVCPort_io_newFlit_x ),
       .io_outPorts_4_x( switch_io_outPorts_4_x ),
       .io_outPorts_3_x( switch_io_outPorts_3_x ),
       .io_outPorts_2_x( switch_io_outPorts_2_x ),
       .io_outPorts_1_x( switch_io_outPorts_1_x ),
       .io_outPorts_0_x( switch_io_outPorts_0_x ),
       .io_sel_4( swAllocator_io_chosens_4 ),
       .io_sel_3( swAllocator_io_chosens_3 ),
       .io_sel_2( swAllocator_io_chosens_2 ),
       .io_sel_1( swAllocator_io_chosens_1 ),
       .io_sel_0( swAllocator_io_chosens_0 )
  );
  SwitchAllocator_0 swAllocator(.clk(clk), .reset(reset),
       .io_requests_4_9_releaseLock( T3092 ),
       .io_requests_4_9_grant( swAllocator_io_requests_4_9_grant ),
       .io_requests_4_9_request( T3088 ),
       .io_requests_4_9_priorityLevel( R2801 ),
       .io_requests_4_8_releaseLock( T3085 ),
       .io_requests_4_8_grant( swAllocator_io_requests_4_8_grant ),
       .io_requests_4_8_request( T3081 ),
       .io_requests_4_8_priorityLevel( R2787 ),
       .io_requests_4_7_releaseLock( T3078 ),
       .io_requests_4_7_grant( swAllocator_io_requests_4_7_grant ),
       .io_requests_4_7_request( T3074 ),
       .io_requests_4_7_priorityLevel( R2773 ),
       .io_requests_4_6_releaseLock( T3071 ),
       .io_requests_4_6_grant( swAllocator_io_requests_4_6_grant ),
       .io_requests_4_6_request( T3067 ),
       .io_requests_4_6_priorityLevel( R2759 ),
       .io_requests_4_5_releaseLock( T3064 ),
       .io_requests_4_5_grant( swAllocator_io_requests_4_5_grant ),
       .io_requests_4_5_request( T3060 ),
       .io_requests_4_5_priorityLevel( R2745 ),
       .io_requests_4_4_releaseLock( T3057 ),
       .io_requests_4_4_grant( swAllocator_io_requests_4_4_grant ),
       .io_requests_4_4_request( T3053 ),
       .io_requests_4_4_priorityLevel( R2731 ),
       .io_requests_4_3_releaseLock( T3050 ),
       .io_requests_4_3_grant( swAllocator_io_requests_4_3_grant ),
       .io_requests_4_3_request( T3046 ),
       .io_requests_4_3_priorityLevel( R2717 ),
       .io_requests_4_2_releaseLock( T3043 ),
       .io_requests_4_2_grant( swAllocator_io_requests_4_2_grant ),
       .io_requests_4_2_request( T3039 ),
       .io_requests_4_2_priorityLevel( R2703 ),
       .io_requests_4_1_releaseLock( T3036 ),
       .io_requests_4_1_grant( swAllocator_io_requests_4_1_grant ),
       .io_requests_4_1_request( T3032 ),
       .io_requests_4_1_priorityLevel( R2689 ),
       .io_requests_4_0_releaseLock( T3029 ),
       .io_requests_4_0_grant( swAllocator_io_requests_4_0_grant ),
       .io_requests_4_0_request( T3025 ),
       .io_requests_4_0_priorityLevel( R2675 ),
       .io_requests_3_9_releaseLock( T3022 ),
       .io_requests_3_9_grant( swAllocator_io_requests_3_9_grant ),
       .io_requests_3_9_request( T3018 ),
       .io_requests_3_9_priorityLevel( R2801 ),
       .io_requests_3_8_releaseLock( T3015 ),
       .io_requests_3_8_grant( swAllocator_io_requests_3_8_grant ),
       .io_requests_3_8_request( T3011 ),
       .io_requests_3_8_priorityLevel( R2787 ),
       .io_requests_3_7_releaseLock( T3008 ),
       .io_requests_3_7_grant( swAllocator_io_requests_3_7_grant ),
       .io_requests_3_7_request( T3004 ),
       .io_requests_3_7_priorityLevel( R2773 ),
       .io_requests_3_6_releaseLock( T3001 ),
       .io_requests_3_6_grant( swAllocator_io_requests_3_6_grant ),
       .io_requests_3_6_request( T2997 ),
       .io_requests_3_6_priorityLevel( R2759 ),
       .io_requests_3_5_releaseLock( T2994 ),
       .io_requests_3_5_grant( swAllocator_io_requests_3_5_grant ),
       .io_requests_3_5_request( T2990 ),
       .io_requests_3_5_priorityLevel( R2745 ),
       .io_requests_3_4_releaseLock( T2987 ),
       .io_requests_3_4_grant( swAllocator_io_requests_3_4_grant ),
       .io_requests_3_4_request( T2983 ),
       .io_requests_3_4_priorityLevel( R2731 ),
       .io_requests_3_3_releaseLock( T2980 ),
       .io_requests_3_3_grant( swAllocator_io_requests_3_3_grant ),
       .io_requests_3_3_request( T2976 ),
       .io_requests_3_3_priorityLevel( R2717 ),
       .io_requests_3_2_releaseLock( T2973 ),
       .io_requests_3_2_grant( swAllocator_io_requests_3_2_grant ),
       .io_requests_3_2_request( T2969 ),
       .io_requests_3_2_priorityLevel( R2703 ),
       .io_requests_3_1_releaseLock( T2966 ),
       .io_requests_3_1_grant( swAllocator_io_requests_3_1_grant ),
       .io_requests_3_1_request( T2962 ),
       .io_requests_3_1_priorityLevel( R2689 ),
       .io_requests_3_0_releaseLock( T2959 ),
       .io_requests_3_0_grant( swAllocator_io_requests_3_0_grant ),
       .io_requests_3_0_request( T2955 ),
       .io_requests_3_0_priorityLevel( R2675 ),
       .io_requests_2_9_releaseLock( T2952 ),
       .io_requests_2_9_grant( swAllocator_io_requests_2_9_grant ),
       .io_requests_2_9_request( T2948 ),
       .io_requests_2_9_priorityLevel( R2801 ),
       .io_requests_2_8_releaseLock( T2945 ),
       .io_requests_2_8_grant( swAllocator_io_requests_2_8_grant ),
       .io_requests_2_8_request( T2941 ),
       .io_requests_2_8_priorityLevel( R2787 ),
       .io_requests_2_7_releaseLock( T2938 ),
       .io_requests_2_7_grant( swAllocator_io_requests_2_7_grant ),
       .io_requests_2_7_request( T2934 ),
       .io_requests_2_7_priorityLevel( R2773 ),
       .io_requests_2_6_releaseLock( T2931 ),
       .io_requests_2_6_grant( swAllocator_io_requests_2_6_grant ),
       .io_requests_2_6_request( T2927 ),
       .io_requests_2_6_priorityLevel( R2759 ),
       .io_requests_2_5_releaseLock( T2924 ),
       .io_requests_2_5_grant( swAllocator_io_requests_2_5_grant ),
       .io_requests_2_5_request( T2920 ),
       .io_requests_2_5_priorityLevel( R2745 ),
       .io_requests_2_4_releaseLock( T2917 ),
       .io_requests_2_4_grant( swAllocator_io_requests_2_4_grant ),
       .io_requests_2_4_request( T2913 ),
       .io_requests_2_4_priorityLevel( R2731 ),
       .io_requests_2_3_releaseLock( T2910 ),
       .io_requests_2_3_grant( swAllocator_io_requests_2_3_grant ),
       .io_requests_2_3_request( T2906 ),
       .io_requests_2_3_priorityLevel( R2717 ),
       .io_requests_2_2_releaseLock( T2903 ),
       .io_requests_2_2_grant( swAllocator_io_requests_2_2_grant ),
       .io_requests_2_2_request( T2899 ),
       .io_requests_2_2_priorityLevel( R2703 ),
       .io_requests_2_1_releaseLock( T2896 ),
       .io_requests_2_1_grant( swAllocator_io_requests_2_1_grant ),
       .io_requests_2_1_request( T2892 ),
       .io_requests_2_1_priorityLevel( R2689 ),
       .io_requests_2_0_releaseLock( T2889 ),
       .io_requests_2_0_grant( swAllocator_io_requests_2_0_grant ),
       .io_requests_2_0_request( T2885 ),
       .io_requests_2_0_priorityLevel( R2675 ),
       .io_requests_1_9_releaseLock( T2882 ),
       .io_requests_1_9_grant( swAllocator_io_requests_1_9_grant ),
       .io_requests_1_9_request( T2878 ),
       .io_requests_1_9_priorityLevel( R2801 ),
       .io_requests_1_8_releaseLock( T2875 ),
       .io_requests_1_8_grant( swAllocator_io_requests_1_8_grant ),
       .io_requests_1_8_request( T2871 ),
       .io_requests_1_8_priorityLevel( R2787 ),
       .io_requests_1_7_releaseLock( T2868 ),
       .io_requests_1_7_grant( swAllocator_io_requests_1_7_grant ),
       .io_requests_1_7_request( T2864 ),
       .io_requests_1_7_priorityLevel( R2773 ),
       .io_requests_1_6_releaseLock( T2861 ),
       .io_requests_1_6_grant( swAllocator_io_requests_1_6_grant ),
       .io_requests_1_6_request( T2857 ),
       .io_requests_1_6_priorityLevel( R2759 ),
       .io_requests_1_5_releaseLock( T2854 ),
       .io_requests_1_5_grant( swAllocator_io_requests_1_5_grant ),
       .io_requests_1_5_request( T2850 ),
       .io_requests_1_5_priorityLevel( R2745 ),
       .io_requests_1_4_releaseLock( T2847 ),
       .io_requests_1_4_grant( swAllocator_io_requests_1_4_grant ),
       .io_requests_1_4_request( T2843 ),
       .io_requests_1_4_priorityLevel( R2731 ),
       .io_requests_1_3_releaseLock( T2840 ),
       .io_requests_1_3_grant( swAllocator_io_requests_1_3_grant ),
       .io_requests_1_3_request( T2836 ),
       .io_requests_1_3_priorityLevel( R2717 ),
       .io_requests_1_2_releaseLock( T2833 ),
       .io_requests_1_2_grant( swAllocator_io_requests_1_2_grant ),
       .io_requests_1_2_request( T2829 ),
       .io_requests_1_2_priorityLevel( R2703 ),
       .io_requests_1_1_releaseLock( T2826 ),
       .io_requests_1_1_grant( swAllocator_io_requests_1_1_grant ),
       .io_requests_1_1_request( T2822 ),
       .io_requests_1_1_priorityLevel( R2689 ),
       .io_requests_1_0_releaseLock( T2819 ),
       .io_requests_1_0_grant( swAllocator_io_requests_1_0_grant ),
       .io_requests_1_0_request( T2815 ),
       .io_requests_1_0_priorityLevel( R2675 ),
       .io_requests_0_9_releaseLock( T2811 ),
       .io_requests_0_9_grant( swAllocator_io_requests_0_9_grant ),
       .io_requests_0_9_request( T2805 ),
       .io_requests_0_9_priorityLevel( R2801 ),
       .io_requests_0_8_releaseLock( T2797 ),
       .io_requests_0_8_grant( swAllocator_io_requests_0_8_grant ),
       .io_requests_0_8_request( T2791 ),
       .io_requests_0_8_priorityLevel( R2787 ),
       .io_requests_0_7_releaseLock( T2783 ),
       .io_requests_0_7_grant( swAllocator_io_requests_0_7_grant ),
       .io_requests_0_7_request( T2777 ),
       .io_requests_0_7_priorityLevel( R2773 ),
       .io_requests_0_6_releaseLock( T2769 ),
       .io_requests_0_6_grant( swAllocator_io_requests_0_6_grant ),
       .io_requests_0_6_request( T2763 ),
       .io_requests_0_6_priorityLevel( R2759 ),
       .io_requests_0_5_releaseLock( T2755 ),
       .io_requests_0_5_grant( swAllocator_io_requests_0_5_grant ),
       .io_requests_0_5_request( T2749 ),
       .io_requests_0_5_priorityLevel( R2745 ),
       .io_requests_0_4_releaseLock( T2741 ),
       .io_requests_0_4_grant( swAllocator_io_requests_0_4_grant ),
       .io_requests_0_4_request( T2735 ),
       .io_requests_0_4_priorityLevel( R2731 ),
       .io_requests_0_3_releaseLock( T2727 ),
       .io_requests_0_3_grant( swAllocator_io_requests_0_3_grant ),
       .io_requests_0_3_request( T2721 ),
       .io_requests_0_3_priorityLevel( R2717 ),
       .io_requests_0_2_releaseLock( T2713 ),
       .io_requests_0_2_grant( swAllocator_io_requests_0_2_grant ),
       .io_requests_0_2_request( T2707 ),
       .io_requests_0_2_priorityLevel( R2703 ),
       .io_requests_0_1_releaseLock( T2699 ),
       .io_requests_0_1_grant( swAllocator_io_requests_0_1_grant ),
       .io_requests_0_1_request( T2693 ),
       .io_requests_0_1_priorityLevel( R2689 ),
       .io_requests_0_0_releaseLock( T2685 ),
       .io_requests_0_0_grant( swAllocator_io_requests_0_0_grant ),
       .io_requests_0_0_request( T2679 ),
       .io_requests_0_0_priorityLevel( R2675 ),
       .io_resources_4_ready( 1'h1 ),
       //.io_resources_4_valid(  )
       .io_resources_3_ready( 1'h1 ),
       //.io_resources_3_valid(  )
       .io_resources_2_ready( 1'h1 ),
       //.io_resources_2_valid(  )
       .io_resources_1_ready( 1'h1 ),
       //.io_resources_1_valid(  )
       .io_resources_0_ready( 1'h1 ),
       //.io_resources_0_valid(  )
       .io_chosens_4( swAllocator_io_chosens_4 ),
       .io_chosens_3( swAllocator_io_chosens_3 ),
       .io_chosens_2( swAllocator_io_chosens_2 ),
       .io_chosens_1( swAllocator_io_chosens_1 ),
       .io_chosens_0( swAllocator_io_chosens_0 )
  );
  SwitchAllocator_1 vcAllocator(.clk(clk), .reset(reset),
       .io_requests_9_9_releaseLock( R2671 ),
       //.io_requests_9_9_grant(  )
       .io_requests_9_9_request( T2670 ),
       //.io_requests_9_9_priorityLevel(  )
       .io_requests_9_8_releaseLock( R2666 ),
       //.io_requests_9_8_grant(  )
       .io_requests_9_8_request( T2665 ),
       //.io_requests_9_8_priorityLevel(  )
       .io_requests_9_7_releaseLock( R2661 ),
       //.io_requests_9_7_grant(  )
       .io_requests_9_7_request( T2660 ),
       //.io_requests_9_7_priorityLevel(  )
       .io_requests_9_6_releaseLock( R2656 ),
       //.io_requests_9_6_grant(  )
       .io_requests_9_6_request( T2655 ),
       //.io_requests_9_6_priorityLevel(  )
       .io_requests_9_5_releaseLock( R2651 ),
       //.io_requests_9_5_grant(  )
       .io_requests_9_5_request( T2650 ),
       //.io_requests_9_5_priorityLevel(  )
       .io_requests_9_4_releaseLock( R2646 ),
       //.io_requests_9_4_grant(  )
       .io_requests_9_4_request( T2645 ),
       //.io_requests_9_4_priorityLevel(  )
       .io_requests_9_3_releaseLock( R2641 ),
       //.io_requests_9_3_grant(  )
       .io_requests_9_3_request( T2640 ),
       //.io_requests_9_3_priorityLevel(  )
       .io_requests_9_2_releaseLock( R2636 ),
       //.io_requests_9_2_grant(  )
       .io_requests_9_2_request( T2635 ),
       //.io_requests_9_2_priorityLevel(  )
       .io_requests_9_1_releaseLock( R2631 ),
       //.io_requests_9_1_grant(  )
       .io_requests_9_1_request( T2630 ),
       //.io_requests_9_1_priorityLevel(  )
       .io_requests_9_0_releaseLock( R2626 ),
       //.io_requests_9_0_grant(  )
       .io_requests_9_0_request( T2625 ),
       //.io_requests_9_0_priorityLevel(  )
       .io_requests_8_9_releaseLock( R2621 ),
       //.io_requests_8_9_grant(  )
       .io_requests_8_9_request( T2620 ),
       //.io_requests_8_9_priorityLevel(  )
       .io_requests_8_8_releaseLock( R2616 ),
       //.io_requests_8_8_grant(  )
       .io_requests_8_8_request( T2615 ),
       //.io_requests_8_8_priorityLevel(  )
       .io_requests_8_7_releaseLock( R2611 ),
       //.io_requests_8_7_grant(  )
       .io_requests_8_7_request( T2610 ),
       //.io_requests_8_7_priorityLevel(  )
       .io_requests_8_6_releaseLock( R2606 ),
       //.io_requests_8_6_grant(  )
       .io_requests_8_6_request( T2605 ),
       //.io_requests_8_6_priorityLevel(  )
       .io_requests_8_5_releaseLock( R2601 ),
       //.io_requests_8_5_grant(  )
       .io_requests_8_5_request( T2600 ),
       //.io_requests_8_5_priorityLevel(  )
       .io_requests_8_4_releaseLock( R2596 ),
       //.io_requests_8_4_grant(  )
       .io_requests_8_4_request( T2595 ),
       //.io_requests_8_4_priorityLevel(  )
       .io_requests_8_3_releaseLock( R2591 ),
       //.io_requests_8_3_grant(  )
       .io_requests_8_3_request( T2590 ),
       //.io_requests_8_3_priorityLevel(  )
       .io_requests_8_2_releaseLock( R2586 ),
       //.io_requests_8_2_grant(  )
       .io_requests_8_2_request( T2585 ),
       //.io_requests_8_2_priorityLevel(  )
       .io_requests_8_1_releaseLock( R2581 ),
       //.io_requests_8_1_grant(  )
       .io_requests_8_1_request( T2580 ),
       //.io_requests_8_1_priorityLevel(  )
       .io_requests_8_0_releaseLock( R2576 ),
       //.io_requests_8_0_grant(  )
       .io_requests_8_0_request( T2575 ),
       //.io_requests_8_0_priorityLevel(  )
       .io_requests_7_9_releaseLock( R2571 ),
       //.io_requests_7_9_grant(  )
       .io_requests_7_9_request( T2570 ),
       //.io_requests_7_9_priorityLevel(  )
       .io_requests_7_8_releaseLock( R2566 ),
       //.io_requests_7_8_grant(  )
       .io_requests_7_8_request( T2565 ),
       //.io_requests_7_8_priorityLevel(  )
       .io_requests_7_7_releaseLock( R2561 ),
       //.io_requests_7_7_grant(  )
       .io_requests_7_7_request( T2560 ),
       //.io_requests_7_7_priorityLevel(  )
       .io_requests_7_6_releaseLock( R2556 ),
       //.io_requests_7_6_grant(  )
       .io_requests_7_6_request( T2555 ),
       //.io_requests_7_6_priorityLevel(  )
       .io_requests_7_5_releaseLock( R2551 ),
       //.io_requests_7_5_grant(  )
       .io_requests_7_5_request( T2550 ),
       //.io_requests_7_5_priorityLevel(  )
       .io_requests_7_4_releaseLock( R2546 ),
       //.io_requests_7_4_grant(  )
       .io_requests_7_4_request( T2545 ),
       //.io_requests_7_4_priorityLevel(  )
       .io_requests_7_3_releaseLock( R2541 ),
       //.io_requests_7_3_grant(  )
       .io_requests_7_3_request( T2540 ),
       //.io_requests_7_3_priorityLevel(  )
       .io_requests_7_2_releaseLock( R2536 ),
       //.io_requests_7_2_grant(  )
       .io_requests_7_2_request( T2535 ),
       //.io_requests_7_2_priorityLevel(  )
       .io_requests_7_1_releaseLock( R2531 ),
       //.io_requests_7_1_grant(  )
       .io_requests_7_1_request( T2530 ),
       //.io_requests_7_1_priorityLevel(  )
       .io_requests_7_0_releaseLock( R2526 ),
       //.io_requests_7_0_grant(  )
       .io_requests_7_0_request( T2525 ),
       //.io_requests_7_0_priorityLevel(  )
       .io_requests_6_9_releaseLock( R2521 ),
       //.io_requests_6_9_grant(  )
       .io_requests_6_9_request( T2520 ),
       //.io_requests_6_9_priorityLevel(  )
       .io_requests_6_8_releaseLock( R2516 ),
       //.io_requests_6_8_grant(  )
       .io_requests_6_8_request( T2515 ),
       //.io_requests_6_8_priorityLevel(  )
       .io_requests_6_7_releaseLock( R2511 ),
       //.io_requests_6_7_grant(  )
       .io_requests_6_7_request( T2510 ),
       //.io_requests_6_7_priorityLevel(  )
       .io_requests_6_6_releaseLock( R2506 ),
       //.io_requests_6_6_grant(  )
       .io_requests_6_6_request( T2505 ),
       //.io_requests_6_6_priorityLevel(  )
       .io_requests_6_5_releaseLock( R2501 ),
       //.io_requests_6_5_grant(  )
       .io_requests_6_5_request( T2500 ),
       //.io_requests_6_5_priorityLevel(  )
       .io_requests_6_4_releaseLock( R2496 ),
       //.io_requests_6_4_grant(  )
       .io_requests_6_4_request( T2495 ),
       //.io_requests_6_4_priorityLevel(  )
       .io_requests_6_3_releaseLock( R2491 ),
       //.io_requests_6_3_grant(  )
       .io_requests_6_3_request( T2490 ),
       //.io_requests_6_3_priorityLevel(  )
       .io_requests_6_2_releaseLock( R2486 ),
       //.io_requests_6_2_grant(  )
       .io_requests_6_2_request( T2485 ),
       //.io_requests_6_2_priorityLevel(  )
       .io_requests_6_1_releaseLock( R2481 ),
       //.io_requests_6_1_grant(  )
       .io_requests_6_1_request( T2480 ),
       //.io_requests_6_1_priorityLevel(  )
       .io_requests_6_0_releaseLock( R2476 ),
       //.io_requests_6_0_grant(  )
       .io_requests_6_0_request( T2475 ),
       //.io_requests_6_0_priorityLevel(  )
       .io_requests_5_9_releaseLock( R2471 ),
       //.io_requests_5_9_grant(  )
       .io_requests_5_9_request( T2470 ),
       //.io_requests_5_9_priorityLevel(  )
       .io_requests_5_8_releaseLock( R2466 ),
       //.io_requests_5_8_grant(  )
       .io_requests_5_8_request( T2465 ),
       //.io_requests_5_8_priorityLevel(  )
       .io_requests_5_7_releaseLock( R2461 ),
       //.io_requests_5_7_grant(  )
       .io_requests_5_7_request( T2460 ),
       //.io_requests_5_7_priorityLevel(  )
       .io_requests_5_6_releaseLock( R2456 ),
       //.io_requests_5_6_grant(  )
       .io_requests_5_6_request( T2455 ),
       //.io_requests_5_6_priorityLevel(  )
       .io_requests_5_5_releaseLock( R2451 ),
       //.io_requests_5_5_grant(  )
       .io_requests_5_5_request( T2450 ),
       //.io_requests_5_5_priorityLevel(  )
       .io_requests_5_4_releaseLock( R2446 ),
       //.io_requests_5_4_grant(  )
       .io_requests_5_4_request( T2445 ),
       //.io_requests_5_4_priorityLevel(  )
       .io_requests_5_3_releaseLock( R2441 ),
       //.io_requests_5_3_grant(  )
       .io_requests_5_3_request( T2440 ),
       //.io_requests_5_3_priorityLevel(  )
       .io_requests_5_2_releaseLock( R2436 ),
       //.io_requests_5_2_grant(  )
       .io_requests_5_2_request( T2435 ),
       //.io_requests_5_2_priorityLevel(  )
       .io_requests_5_1_releaseLock( R2431 ),
       //.io_requests_5_1_grant(  )
       .io_requests_5_1_request( T2430 ),
       //.io_requests_5_1_priorityLevel(  )
       .io_requests_5_0_releaseLock( R2426 ),
       //.io_requests_5_0_grant(  )
       .io_requests_5_0_request( T2425 ),
       //.io_requests_5_0_priorityLevel(  )
       .io_requests_4_9_releaseLock( R2421 ),
       //.io_requests_4_9_grant(  )
       .io_requests_4_9_request( T2420 ),
       //.io_requests_4_9_priorityLevel(  )
       .io_requests_4_8_releaseLock( R2416 ),
       //.io_requests_4_8_grant(  )
       .io_requests_4_8_request( T2415 ),
       //.io_requests_4_8_priorityLevel(  )
       .io_requests_4_7_releaseLock( R2411 ),
       //.io_requests_4_7_grant(  )
       .io_requests_4_7_request( T2410 ),
       //.io_requests_4_7_priorityLevel(  )
       .io_requests_4_6_releaseLock( R2406 ),
       //.io_requests_4_6_grant(  )
       .io_requests_4_6_request( T2405 ),
       //.io_requests_4_6_priorityLevel(  )
       .io_requests_4_5_releaseLock( R2401 ),
       //.io_requests_4_5_grant(  )
       .io_requests_4_5_request( T2400 ),
       //.io_requests_4_5_priorityLevel(  )
       .io_requests_4_4_releaseLock( R2396 ),
       //.io_requests_4_4_grant(  )
       .io_requests_4_4_request( T2395 ),
       //.io_requests_4_4_priorityLevel(  )
       .io_requests_4_3_releaseLock( R2391 ),
       //.io_requests_4_3_grant(  )
       .io_requests_4_3_request( T2390 ),
       //.io_requests_4_3_priorityLevel(  )
       .io_requests_4_2_releaseLock( R2386 ),
       //.io_requests_4_2_grant(  )
       .io_requests_4_2_request( T2385 ),
       //.io_requests_4_2_priorityLevel(  )
       .io_requests_4_1_releaseLock( R2381 ),
       //.io_requests_4_1_grant(  )
       .io_requests_4_1_request( T2380 ),
       //.io_requests_4_1_priorityLevel(  )
       .io_requests_4_0_releaseLock( R2376 ),
       //.io_requests_4_0_grant(  )
       .io_requests_4_0_request( T2375 ),
       //.io_requests_4_0_priorityLevel(  )
       .io_requests_3_9_releaseLock( R2371 ),
       //.io_requests_3_9_grant(  )
       .io_requests_3_9_request( T2370 ),
       //.io_requests_3_9_priorityLevel(  )
       .io_requests_3_8_releaseLock( R2366 ),
       //.io_requests_3_8_grant(  )
       .io_requests_3_8_request( T2365 ),
       //.io_requests_3_8_priorityLevel(  )
       .io_requests_3_7_releaseLock( R2361 ),
       //.io_requests_3_7_grant(  )
       .io_requests_3_7_request( T2360 ),
       //.io_requests_3_7_priorityLevel(  )
       .io_requests_3_6_releaseLock( R2356 ),
       //.io_requests_3_6_grant(  )
       .io_requests_3_6_request( T2355 ),
       //.io_requests_3_6_priorityLevel(  )
       .io_requests_3_5_releaseLock( R2351 ),
       //.io_requests_3_5_grant(  )
       .io_requests_3_5_request( T2350 ),
       //.io_requests_3_5_priorityLevel(  )
       .io_requests_3_4_releaseLock( R2346 ),
       //.io_requests_3_4_grant(  )
       .io_requests_3_4_request( T2345 ),
       //.io_requests_3_4_priorityLevel(  )
       .io_requests_3_3_releaseLock( R2341 ),
       //.io_requests_3_3_grant(  )
       .io_requests_3_3_request( T2340 ),
       //.io_requests_3_3_priorityLevel(  )
       .io_requests_3_2_releaseLock( R2336 ),
       //.io_requests_3_2_grant(  )
       .io_requests_3_2_request( T2335 ),
       //.io_requests_3_2_priorityLevel(  )
       .io_requests_3_1_releaseLock( R2331 ),
       //.io_requests_3_1_grant(  )
       .io_requests_3_1_request( T2330 ),
       //.io_requests_3_1_priorityLevel(  )
       .io_requests_3_0_releaseLock( R2326 ),
       //.io_requests_3_0_grant(  )
       .io_requests_3_0_request( T2325 ),
       //.io_requests_3_0_priorityLevel(  )
       .io_requests_2_9_releaseLock( R2321 ),
       //.io_requests_2_9_grant(  )
       .io_requests_2_9_request( T2320 ),
       //.io_requests_2_9_priorityLevel(  )
       .io_requests_2_8_releaseLock( R2316 ),
       //.io_requests_2_8_grant(  )
       .io_requests_2_8_request( T2315 ),
       //.io_requests_2_8_priorityLevel(  )
       .io_requests_2_7_releaseLock( R2311 ),
       //.io_requests_2_7_grant(  )
       .io_requests_2_7_request( T2310 ),
       //.io_requests_2_7_priorityLevel(  )
       .io_requests_2_6_releaseLock( R2306 ),
       //.io_requests_2_6_grant(  )
       .io_requests_2_6_request( T2305 ),
       //.io_requests_2_6_priorityLevel(  )
       .io_requests_2_5_releaseLock( R2301 ),
       //.io_requests_2_5_grant(  )
       .io_requests_2_5_request( T2300 ),
       //.io_requests_2_5_priorityLevel(  )
       .io_requests_2_4_releaseLock( R2296 ),
       //.io_requests_2_4_grant(  )
       .io_requests_2_4_request( T2295 ),
       //.io_requests_2_4_priorityLevel(  )
       .io_requests_2_3_releaseLock( R2291 ),
       //.io_requests_2_3_grant(  )
       .io_requests_2_3_request( T2290 ),
       //.io_requests_2_3_priorityLevel(  )
       .io_requests_2_2_releaseLock( R2286 ),
       //.io_requests_2_2_grant(  )
       .io_requests_2_2_request( T2285 ),
       //.io_requests_2_2_priorityLevel(  )
       .io_requests_2_1_releaseLock( R2281 ),
       //.io_requests_2_1_grant(  )
       .io_requests_2_1_request( T2280 ),
       //.io_requests_2_1_priorityLevel(  )
       .io_requests_2_0_releaseLock( R2276 ),
       //.io_requests_2_0_grant(  )
       .io_requests_2_0_request( T2275 ),
       //.io_requests_2_0_priorityLevel(  )
       .io_requests_1_9_releaseLock( R2271 ),
       //.io_requests_1_9_grant(  )
       .io_requests_1_9_request( T2270 ),
       //.io_requests_1_9_priorityLevel(  )
       .io_requests_1_8_releaseLock( R2266 ),
       //.io_requests_1_8_grant(  )
       .io_requests_1_8_request( T2265 ),
       //.io_requests_1_8_priorityLevel(  )
       .io_requests_1_7_releaseLock( R2261 ),
       //.io_requests_1_7_grant(  )
       .io_requests_1_7_request( T2260 ),
       //.io_requests_1_7_priorityLevel(  )
       .io_requests_1_6_releaseLock( R2256 ),
       //.io_requests_1_6_grant(  )
       .io_requests_1_6_request( T2255 ),
       //.io_requests_1_6_priorityLevel(  )
       .io_requests_1_5_releaseLock( R2251 ),
       //.io_requests_1_5_grant(  )
       .io_requests_1_5_request( T2250 ),
       //.io_requests_1_5_priorityLevel(  )
       .io_requests_1_4_releaseLock( R2246 ),
       //.io_requests_1_4_grant(  )
       .io_requests_1_4_request( T2245 ),
       //.io_requests_1_4_priorityLevel(  )
       .io_requests_1_3_releaseLock( R2241 ),
       //.io_requests_1_3_grant(  )
       .io_requests_1_3_request( T2240 ),
       //.io_requests_1_3_priorityLevel(  )
       .io_requests_1_2_releaseLock( R2236 ),
       //.io_requests_1_2_grant(  )
       .io_requests_1_2_request( T2235 ),
       //.io_requests_1_2_priorityLevel(  )
       .io_requests_1_1_releaseLock( R2231 ),
       //.io_requests_1_1_grant(  )
       .io_requests_1_1_request( T2230 ),
       //.io_requests_1_1_priorityLevel(  )
       .io_requests_1_0_releaseLock( R2226 ),
       //.io_requests_1_0_grant(  )
       .io_requests_1_0_request( T2225 ),
       //.io_requests_1_0_priorityLevel(  )
       .io_requests_0_9_releaseLock( R2221 ),
       //.io_requests_0_9_grant(  )
       .io_requests_0_9_request( T2220 ),
       //.io_requests_0_9_priorityLevel(  )
       .io_requests_0_8_releaseLock( R2216 ),
       //.io_requests_0_8_grant(  )
       .io_requests_0_8_request( T2215 ),
       //.io_requests_0_8_priorityLevel(  )
       .io_requests_0_7_releaseLock( R2211 ),
       //.io_requests_0_7_grant(  )
       .io_requests_0_7_request( T2210 ),
       //.io_requests_0_7_priorityLevel(  )
       .io_requests_0_6_releaseLock( R2206 ),
       //.io_requests_0_6_grant(  )
       .io_requests_0_6_request( T2205 ),
       //.io_requests_0_6_priorityLevel(  )
       .io_requests_0_5_releaseLock( R2201 ),
       //.io_requests_0_5_grant(  )
       .io_requests_0_5_request( T2200 ),
       //.io_requests_0_5_priorityLevel(  )
       .io_requests_0_4_releaseLock( R2196 ),
       //.io_requests_0_4_grant(  )
       .io_requests_0_4_request( T2195 ),
       //.io_requests_0_4_priorityLevel(  )
       .io_requests_0_3_releaseLock( R2191 ),
       //.io_requests_0_3_grant(  )
       .io_requests_0_3_request( T2190 ),
       //.io_requests_0_3_priorityLevel(  )
       .io_requests_0_2_releaseLock( R2186 ),
       //.io_requests_0_2_grant(  )
       .io_requests_0_2_request( T2185 ),
       //.io_requests_0_2_priorityLevel(  )
       .io_requests_0_1_releaseLock( R2181 ),
       //.io_requests_0_1_grant(  )
       .io_requests_0_1_request( T2180 ),
       //.io_requests_0_1_priorityLevel(  )
       .io_requests_0_0_releaseLock( R2176 ),
       //.io_requests_0_0_grant(  )
       .io_requests_0_0_request( T2175 ),
       //.io_requests_0_0_priorityLevel(  )
       .io_resources_9_ready( T2173 ),
       .io_resources_9_valid( vcAllocator_io_resources_9_valid ),
       .io_resources_8_ready( T2171 ),
       .io_resources_8_valid( vcAllocator_io_resources_8_valid ),
       .io_resources_7_ready( T2169 ),
       .io_resources_7_valid( vcAllocator_io_resources_7_valid ),
       .io_resources_6_ready( T2167 ),
       .io_resources_6_valid( vcAllocator_io_resources_6_valid ),
       .io_resources_5_ready( T2165 ),
       .io_resources_5_valid( vcAllocator_io_resources_5_valid ),
       .io_resources_4_ready( T2163 ),
       .io_resources_4_valid( vcAllocator_io_resources_4_valid ),
       .io_resources_3_ready( T2161 ),
       .io_resources_3_valid( vcAllocator_io_resources_3_valid ),
       .io_resources_2_ready( T2159 ),
       .io_resources_2_valid( vcAllocator_io_resources_2_valid ),
       .io_resources_1_ready( T2157 ),
       .io_resources_1_valid( vcAllocator_io_resources_1_valid ),
       .io_resources_0_ready( T2155 ),
       .io_resources_0_valid( vcAllocator_io_resources_0_valid ),
       .io_chosens_9( vcAllocator_io_chosens_9 ),
       .io_chosens_8( vcAllocator_io_chosens_8 ),
       .io_chosens_7( vcAllocator_io_chosens_7 ),
       .io_chosens_6( vcAllocator_io_chosens_6 ),
       .io_chosens_5( vcAllocator_io_chosens_5 ),
       .io_chosens_4( vcAllocator_io_chosens_4 ),
       .io_chosens_3( vcAllocator_io_chosens_3 ),
       .io_chosens_2( vcAllocator_io_chosens_2 ),
       .io_chosens_1( vcAllocator_io_chosens_1 ),
       .io_chosens_0( vcAllocator_io_chosens_0 )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign vcAllocator.io_requests_9_9_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_9_8_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_9_7_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_9_6_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_9_5_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_9_4_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_9_3_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_9_2_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_9_1_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_9_0_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_8_9_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_8_8_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_8_7_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_8_6_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_8_5_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_8_4_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_8_3_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_8_2_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_8_1_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_8_0_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_7_9_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_7_8_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_7_7_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_7_6_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_7_5_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_7_4_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_7_3_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_7_2_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_7_1_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_7_0_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_6_9_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_6_8_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_6_7_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_6_6_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_6_5_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_6_4_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_6_3_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_6_2_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_6_1_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_6_0_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_5_9_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_5_8_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_5_7_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_5_6_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_5_5_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_5_4_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_5_3_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_5_2_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_5_1_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_5_0_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_4_9_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_4_8_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_4_7_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_4_6_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_4_5_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_4_4_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_4_3_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_4_2_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_4_1_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_4_0_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_3_9_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_3_8_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_3_7_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_3_6_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_3_5_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_3_4_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_3_3_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_3_2_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_3_1_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_3_0_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_2_9_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_2_8_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_2_7_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_2_6_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_2_5_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_2_4_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_2_3_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_2_2_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_2_1_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_2_0_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_1_9_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_1_8_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_1_7_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_1_6_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_1_5_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_1_4_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_1_3_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_1_2_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_1_1_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_1_0_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_0_9_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_0_8_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_0_7_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_0_6_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_0_5_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_0_4_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_0_3_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_0_2_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_0_1_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_0_0_priorityLevel = {1{1'b0}};
// synthesis translate_on
`endif
  VCRouterOutputStateManagement VCRouterOutputStateManagement(.clk(clk), .reset(reset),
       .io_swAllocGranted( T2094 ),
       .io_creditsAvail( T2092 ),
       .io_currentState( VCRouterOutputStateManagement_io_currentState )
  );
  VCRouterOutputStateManagement VCRouterOutputStateManagement_1(.clk(clk), .reset(reset),
       .io_swAllocGranted( T2031 ),
       .io_creditsAvail( T2029 ),
       .io_currentState( VCRouterOutputStateManagement_1_io_currentState )
  );
  VCRouterOutputStateManagement VCRouterOutputStateManagement_2(.clk(clk), .reset(reset),
       .io_swAllocGranted( T1968 ),
       .io_creditsAvail( T1966 ),
       .io_currentState( VCRouterOutputStateManagement_2_io_currentState )
  );
  VCRouterOutputStateManagement VCRouterOutputStateManagement_3(.clk(clk), .reset(reset),
       .io_swAllocGranted( T1905 ),
       .io_creditsAvail( T1903 ),
       .io_currentState( VCRouterOutputStateManagement_3_io_currentState )
  );
  VCRouterOutputStateManagement VCRouterOutputStateManagement_4(.clk(clk), .reset(reset),
       .io_swAllocGranted( T1722 ),
       .io_creditsAvail( T1720 ),
       .io_currentState( VCRouterOutputStateManagement_4_io_currentState )
  );
  CreditGen CreditGen(
       .io_outCredit_grant( CreditGen_io_outCredit_grant ),
       .io_inGrant( T1710 )
  );
  RouterRegFile RouterRegFile(.clk(clk), .reset(reset),
       .io_writeData( T1708 ),
       .io_writeEnable( T1705 ),
       //.io_full(  )
       .io_readData( RouterRegFile_io_readData ),
       .io_readValid( RouterRegFile_io_readValid ),
       .io_readIncrement( T1692 ),
       .io_writePipelineReg_2( RouterRegFile_io_readPipelineReg_1 ),
       .io_writePipelineReg_1( RouterRegFile_io_readPipelineReg_0 ),
       .io_writePipelineReg_0( T3181 ),
       .io_wePipelineReg_2( T1681 ),
       .io_wePipelineReg_1( T1678 ),
       .io_wePipelineReg_0( T1676 ),
       //.io_readPipelineReg_2(  )
       .io_readPipelineReg_1( RouterRegFile_io_readPipelineReg_1 ),
       .io_readPipelineReg_0( RouterRegFile_io_readPipelineReg_0 ),
       //.io_rvPipelineReg_2(  )
       .io_rvPipelineReg_1( RouterRegFile_io_rvPipelineReg_1 ),
       .io_rvPipelineReg_0( RouterRegFile_io_rvPipelineReg_0 )
  );
  RouterBuffer RouterBuffer(.clk(clk), .reset(reset),
       .io_enq_ready( RouterBuffer_io_enq_ready ),
       .io_enq_valid( T1675 ),
       .io_enq_bits_x( io_inChannels_0_flit_x ),
       .io_deq_ready( T1656 ),
       .io_deq_valid( RouterBuffer_io_deq_valid ),
       .io_deq_bits_x( RouterBuffer_io_deq_bits_x )
  );
  CMeshDOR_0 CMeshDOR(
       .io_inHeadFlit_packetID( T1655 ),
       .io_inHeadFlit_isTail( T1654 ),
       .io_inHeadFlit_vcPort( T1653 ),
       .io_inHeadFlit_packetType( T1652 ),
       .io_inHeadFlit_destination_2( T1651 ),
       .io_inHeadFlit_destination_1( T1650 ),
       .io_inHeadFlit_destination_0( T1649 ),
       .io_inHeadFlit_priorityLevel( T1646 ),
       .io_outHeadFlit_packetID( CMeshDOR_io_outHeadFlit_packetID ),
       .io_outHeadFlit_isTail( CMeshDOR_io_outHeadFlit_isTail ),
       .io_outHeadFlit_vcPort( CMeshDOR_io_outHeadFlit_vcPort ),
       .io_outHeadFlit_packetType( CMeshDOR_io_outHeadFlit_packetType ),
       .io_outHeadFlit_destination_2( CMeshDOR_io_outHeadFlit_destination_2 ),
       .io_outHeadFlit_destination_1( CMeshDOR_io_outHeadFlit_destination_1 ),
       .io_outHeadFlit_destination_0( CMeshDOR_io_outHeadFlit_destination_0 ),
       .io_outHeadFlit_priorityLevel( CMeshDOR_io_outHeadFlit_priorityLevel ),
       .io_result( CMeshDOR_io_result ),
       .io_vcsAvailable_4( CMeshDOR_io_vcsAvailable_4 ),
       .io_vcsAvailable_3( CMeshDOR_io_vcsAvailable_3 ),
       .io_vcsAvailable_2( CMeshDOR_io_vcsAvailable_2 ),
       .io_vcsAvailable_1( CMeshDOR_io_vcsAvailable_1 ),
       .io_vcsAvailable_0( CMeshDOR_io_vcsAvailable_0 )
  );
  VCRouterStateManagement VCRouterStateManagement(.clk(clk), .reset(reset),
       .io_inputBufferValid( RouterBuffer_io_deq_valid ),
       .io_routingComplete( R1645 ),
       .io_inputBufferIsTail( T1636 ),
       .io_vcAllocGranted( vcAllocator_io_resources_0_valid ),
       .io_swAllocGranted( T1616 ),
       .io_creditsAvail( T1597 ),
       .io_outputReady( T1584 ),
       .io_currentState( VCRouterStateManagement_io_currentState )
  );
  ReplaceVCPort ReplaceVCPort(
       .io_oldFlit_x( T1582 ),
       .io_newVCPort( T3175 ),
       .io_newFlit_x( ReplaceVCPort_io_newFlit_x )
  );
  Flit2FlitBundle Flit2FlitBundle(
       .io_inFlit_x( T1576 )
       //.io_outHead_packetID(  )
       //.io_outHead_isTail(  )
       //.io_outHead_vcPort(  )
       //.io_outHead_packetType(  )
       //.io_outHead_destination_2(  )
       //.io_outHead_destination_1(  )
       //.io_outHead_destination_0(  )
       //.io_outHead_priorityLevel(  )
       //.io_outBody_packetID(  )
       //.io_outBody_isTail(  )
       //.io_outBody_vcPort(  )
       //.io_outBody_flitID(  )
       //.io_outBody_payload(  )
  );
  CreditGen CreditGen_1(
       .io_outCredit_grant( CreditGen_1_io_outCredit_grant ),
       .io_inGrant( T1566 )
  );
  RouterRegFile RouterRegFile_1(.clk(clk), .reset(reset),
       .io_writeData( T1564 ),
       .io_writeEnable( T1561 ),
       //.io_full(  )
       .io_readData( RouterRegFile_1_io_readData ),
       .io_readValid( RouterRegFile_1_io_readValid ),
       .io_readIncrement( T1548 ),
       .io_writePipelineReg_2( RouterRegFile_1_io_readPipelineReg_1 ),
       .io_writePipelineReg_1( RouterRegFile_1_io_readPipelineReg_0 ),
       .io_writePipelineReg_0( T3174 ),
       .io_wePipelineReg_2( T1537 ),
       .io_wePipelineReg_1( T1534 ),
       .io_wePipelineReg_0( T1532 ),
       //.io_readPipelineReg_2(  )
       .io_readPipelineReg_1( RouterRegFile_1_io_readPipelineReg_1 ),
       .io_readPipelineReg_0( RouterRegFile_1_io_readPipelineReg_0 ),
       //.io_rvPipelineReg_2(  )
       .io_rvPipelineReg_1( RouterRegFile_1_io_rvPipelineReg_1 ),
       .io_rvPipelineReg_0( RouterRegFile_1_io_rvPipelineReg_0 )
  );
  RouterBuffer RouterBuffer_1(.clk(clk), .reset(reset),
       .io_enq_ready( RouterBuffer_1_io_enq_ready ),
       .io_enq_valid( T1531 ),
       .io_enq_bits_x( io_inChannels_0_flit_x ),
       .io_deq_ready( T1512 ),
       .io_deq_valid( RouterBuffer_1_io_deq_valid ),
       .io_deq_bits_x( RouterBuffer_1_io_deq_bits_x )
  );
  CMeshDOR_0 CMeshDOR_1(
       .io_inHeadFlit_packetID( T1511 ),
       .io_inHeadFlit_isTail( T1510 ),
       .io_inHeadFlit_vcPort( T1509 ),
       .io_inHeadFlit_packetType( T1508 ),
       .io_inHeadFlit_destination_2( T1507 ),
       .io_inHeadFlit_destination_1( T1506 ),
       .io_inHeadFlit_destination_0( T1505 ),
       .io_inHeadFlit_priorityLevel( T1502 ),
       .io_outHeadFlit_packetID( CMeshDOR_1_io_outHeadFlit_packetID ),
       .io_outHeadFlit_isTail( CMeshDOR_1_io_outHeadFlit_isTail ),
       .io_outHeadFlit_vcPort( CMeshDOR_1_io_outHeadFlit_vcPort ),
       .io_outHeadFlit_packetType( CMeshDOR_1_io_outHeadFlit_packetType ),
       .io_outHeadFlit_destination_2( CMeshDOR_1_io_outHeadFlit_destination_2 ),
       .io_outHeadFlit_destination_1( CMeshDOR_1_io_outHeadFlit_destination_1 ),
       .io_outHeadFlit_destination_0( CMeshDOR_1_io_outHeadFlit_destination_0 ),
       .io_outHeadFlit_priorityLevel( CMeshDOR_1_io_outHeadFlit_priorityLevel ),
       .io_result( CMeshDOR_1_io_result ),
       .io_vcsAvailable_4( CMeshDOR_1_io_vcsAvailable_4 ),
       .io_vcsAvailable_3( CMeshDOR_1_io_vcsAvailable_3 ),
       .io_vcsAvailable_2( CMeshDOR_1_io_vcsAvailable_2 ),
       .io_vcsAvailable_1( CMeshDOR_1_io_vcsAvailable_1 ),
       .io_vcsAvailable_0( CMeshDOR_1_io_vcsAvailable_0 )
  );
  VCRouterStateManagement VCRouterStateManagement_1(.clk(clk), .reset(reset),
       .io_inputBufferValid( RouterBuffer_1_io_deq_valid ),
       .io_routingComplete( R1501 ),
       .io_inputBufferIsTail( T1492 ),
       .io_vcAllocGranted( vcAllocator_io_resources_1_valid ),
       .io_swAllocGranted( T1472 ),
       .io_creditsAvail( T1453 ),
       .io_outputReady( T1440 ),
       .io_currentState( VCRouterStateManagement_1_io_currentState )
  );
  ReplaceVCPort ReplaceVCPort_1(
       .io_oldFlit_x( T1438 ),
       .io_newVCPort( T3168 ),
       .io_newFlit_x( ReplaceVCPort_1_io_newFlit_x )
  );
  Flit2FlitBundle Flit2FlitBundle_1(
       .io_inFlit_x( T1432 )
       //.io_outHead_packetID(  )
       //.io_outHead_isTail(  )
       //.io_outHead_vcPort(  )
       //.io_outHead_packetType(  )
       //.io_outHead_destination_2(  )
       //.io_outHead_destination_1(  )
       //.io_outHead_destination_0(  )
       //.io_outHead_priorityLevel(  )
       //.io_outBody_packetID(  )
       //.io_outBody_isTail(  )
       //.io_outBody_vcPort(  )
       //.io_outBody_flitID(  )
       //.io_outBody_payload(  )
  );
  CreditGen CreditGen_2(
       .io_outCredit_grant( CreditGen_2_io_outCredit_grant ),
       .io_inGrant( T1422 )
  );
  RouterRegFile RouterRegFile_2(.clk(clk), .reset(reset),
       .io_writeData( T1420 ),
       .io_writeEnable( T1417 ),
       //.io_full(  )
       .io_readData( RouterRegFile_2_io_readData ),
       .io_readValid( RouterRegFile_2_io_readValid ),
       .io_readIncrement( T1404 ),
       .io_writePipelineReg_2( RouterRegFile_2_io_readPipelineReg_1 ),
       .io_writePipelineReg_1( RouterRegFile_2_io_readPipelineReg_0 ),
       .io_writePipelineReg_0( T3167 ),
       .io_wePipelineReg_2( T1393 ),
       .io_wePipelineReg_1( T1390 ),
       .io_wePipelineReg_0( T1388 ),
       //.io_readPipelineReg_2(  )
       .io_readPipelineReg_1( RouterRegFile_2_io_readPipelineReg_1 ),
       .io_readPipelineReg_0( RouterRegFile_2_io_readPipelineReg_0 ),
       //.io_rvPipelineReg_2(  )
       .io_rvPipelineReg_1( RouterRegFile_2_io_rvPipelineReg_1 ),
       .io_rvPipelineReg_0( RouterRegFile_2_io_rvPipelineReg_0 )
  );
  RouterBuffer RouterBuffer_2(.clk(clk), .reset(reset),
       .io_enq_ready( RouterBuffer_2_io_enq_ready ),
       .io_enq_valid( T1387 ),
       .io_enq_bits_x( io_inChannels_1_flit_x ),
       .io_deq_ready( T1368 ),
       .io_deq_valid( RouterBuffer_2_io_deq_valid ),
       .io_deq_bits_x( RouterBuffer_2_io_deq_bits_x )
  );
  CMeshDOR_0 CMeshDOR_2(
       .io_inHeadFlit_packetID( T1367 ),
       .io_inHeadFlit_isTail( T1366 ),
       .io_inHeadFlit_vcPort( T1365 ),
       .io_inHeadFlit_packetType( T1364 ),
       .io_inHeadFlit_destination_2( T1363 ),
       .io_inHeadFlit_destination_1( T1362 ),
       .io_inHeadFlit_destination_0( T1361 ),
       .io_inHeadFlit_priorityLevel( T1358 ),
       .io_outHeadFlit_packetID( CMeshDOR_2_io_outHeadFlit_packetID ),
       .io_outHeadFlit_isTail( CMeshDOR_2_io_outHeadFlit_isTail ),
       .io_outHeadFlit_vcPort( CMeshDOR_2_io_outHeadFlit_vcPort ),
       .io_outHeadFlit_packetType( CMeshDOR_2_io_outHeadFlit_packetType ),
       .io_outHeadFlit_destination_2( CMeshDOR_2_io_outHeadFlit_destination_2 ),
       .io_outHeadFlit_destination_1( CMeshDOR_2_io_outHeadFlit_destination_1 ),
       .io_outHeadFlit_destination_0( CMeshDOR_2_io_outHeadFlit_destination_0 ),
       .io_outHeadFlit_priorityLevel( CMeshDOR_2_io_outHeadFlit_priorityLevel ),
       .io_result( CMeshDOR_2_io_result ),
       .io_vcsAvailable_4( CMeshDOR_2_io_vcsAvailable_4 ),
       .io_vcsAvailable_3( CMeshDOR_2_io_vcsAvailable_3 ),
       .io_vcsAvailable_2( CMeshDOR_2_io_vcsAvailable_2 ),
       .io_vcsAvailable_1( CMeshDOR_2_io_vcsAvailable_1 ),
       .io_vcsAvailable_0( CMeshDOR_2_io_vcsAvailable_0 )
  );
  VCRouterStateManagement VCRouterStateManagement_2(.clk(clk), .reset(reset),
       .io_inputBufferValid( RouterBuffer_2_io_deq_valid ),
       .io_routingComplete( R1357 ),
       .io_inputBufferIsTail( T1348 ),
       .io_vcAllocGranted( vcAllocator_io_resources_2_valid ),
       .io_swAllocGranted( T1328 ),
       .io_creditsAvail( T1309 ),
       .io_outputReady( T1296 ),
       .io_currentState( VCRouterStateManagement_2_io_currentState )
  );
  ReplaceVCPort ReplaceVCPort_2(
       .io_oldFlit_x( T1294 ),
       .io_newVCPort( T3161 ),
       .io_newFlit_x( ReplaceVCPort_2_io_newFlit_x )
  );
  Flit2FlitBundle Flit2FlitBundle_2(
       .io_inFlit_x( T1288 )
       //.io_outHead_packetID(  )
       //.io_outHead_isTail(  )
       //.io_outHead_vcPort(  )
       //.io_outHead_packetType(  )
       //.io_outHead_destination_2(  )
       //.io_outHead_destination_1(  )
       //.io_outHead_destination_0(  )
       //.io_outHead_priorityLevel(  )
       //.io_outBody_packetID(  )
       //.io_outBody_isTail(  )
       //.io_outBody_vcPort(  )
       //.io_outBody_flitID(  )
       //.io_outBody_payload(  )
  );
  CreditGen CreditGen_3(
       .io_outCredit_grant( CreditGen_3_io_outCredit_grant ),
       .io_inGrant( T1278 )
  );
  RouterRegFile RouterRegFile_3(.clk(clk), .reset(reset),
       .io_writeData( T1276 ),
       .io_writeEnable( T1273 ),
       //.io_full(  )
       .io_readData( RouterRegFile_3_io_readData ),
       .io_readValid( RouterRegFile_3_io_readValid ),
       .io_readIncrement( T1260 ),
       .io_writePipelineReg_2( RouterRegFile_3_io_readPipelineReg_1 ),
       .io_writePipelineReg_1( RouterRegFile_3_io_readPipelineReg_0 ),
       .io_writePipelineReg_0( T3160 ),
       .io_wePipelineReg_2( T1249 ),
       .io_wePipelineReg_1( T1246 ),
       .io_wePipelineReg_0( T1244 ),
       //.io_readPipelineReg_2(  )
       .io_readPipelineReg_1( RouterRegFile_3_io_readPipelineReg_1 ),
       .io_readPipelineReg_0( RouterRegFile_3_io_readPipelineReg_0 ),
       //.io_rvPipelineReg_2(  )
       .io_rvPipelineReg_1( RouterRegFile_3_io_rvPipelineReg_1 ),
       .io_rvPipelineReg_0( RouterRegFile_3_io_rvPipelineReg_0 )
  );
  RouterBuffer RouterBuffer_3(.clk(clk), .reset(reset),
       .io_enq_ready( RouterBuffer_3_io_enq_ready ),
       .io_enq_valid( T1243 ),
       .io_enq_bits_x( io_inChannels_1_flit_x ),
       .io_deq_ready( T1224 ),
       .io_deq_valid( RouterBuffer_3_io_deq_valid ),
       .io_deq_bits_x( RouterBuffer_3_io_deq_bits_x )
  );
  CMeshDOR_0 CMeshDOR_3(
       .io_inHeadFlit_packetID( T1223 ),
       .io_inHeadFlit_isTail( T1222 ),
       .io_inHeadFlit_vcPort( T1221 ),
       .io_inHeadFlit_packetType( T1220 ),
       .io_inHeadFlit_destination_2( T1219 ),
       .io_inHeadFlit_destination_1( T1218 ),
       .io_inHeadFlit_destination_0( T1217 ),
       .io_inHeadFlit_priorityLevel( T1214 ),
       .io_outHeadFlit_packetID( CMeshDOR_3_io_outHeadFlit_packetID ),
       .io_outHeadFlit_isTail( CMeshDOR_3_io_outHeadFlit_isTail ),
       .io_outHeadFlit_vcPort( CMeshDOR_3_io_outHeadFlit_vcPort ),
       .io_outHeadFlit_packetType( CMeshDOR_3_io_outHeadFlit_packetType ),
       .io_outHeadFlit_destination_2( CMeshDOR_3_io_outHeadFlit_destination_2 ),
       .io_outHeadFlit_destination_1( CMeshDOR_3_io_outHeadFlit_destination_1 ),
       .io_outHeadFlit_destination_0( CMeshDOR_3_io_outHeadFlit_destination_0 ),
       .io_outHeadFlit_priorityLevel( CMeshDOR_3_io_outHeadFlit_priorityLevel ),
       .io_result( CMeshDOR_3_io_result ),
       .io_vcsAvailable_4( CMeshDOR_3_io_vcsAvailable_4 ),
       .io_vcsAvailable_3( CMeshDOR_3_io_vcsAvailable_3 ),
       .io_vcsAvailable_2( CMeshDOR_3_io_vcsAvailable_2 ),
       .io_vcsAvailable_1( CMeshDOR_3_io_vcsAvailable_1 ),
       .io_vcsAvailable_0( CMeshDOR_3_io_vcsAvailable_0 )
  );
  VCRouterStateManagement VCRouterStateManagement_3(.clk(clk), .reset(reset),
       .io_inputBufferValid( RouterBuffer_3_io_deq_valid ),
       .io_routingComplete( R1213 ),
       .io_inputBufferIsTail( T1204 ),
       .io_vcAllocGranted( vcAllocator_io_resources_3_valid ),
       .io_swAllocGranted( T1184 ),
       .io_creditsAvail( T1165 ),
       .io_outputReady( T1152 ),
       .io_currentState( VCRouterStateManagement_3_io_currentState )
  );
  ReplaceVCPort ReplaceVCPort_3(
       .io_oldFlit_x( T1150 ),
       .io_newVCPort( T3154 ),
       .io_newFlit_x( ReplaceVCPort_3_io_newFlit_x )
  );
  Flit2FlitBundle Flit2FlitBundle_3(
       .io_inFlit_x( T1144 )
       //.io_outHead_packetID(  )
       //.io_outHead_isTail(  )
       //.io_outHead_vcPort(  )
       //.io_outHead_packetType(  )
       //.io_outHead_destination_2(  )
       //.io_outHead_destination_1(  )
       //.io_outHead_destination_0(  )
       //.io_outHead_priorityLevel(  )
       //.io_outBody_packetID(  )
       //.io_outBody_isTail(  )
       //.io_outBody_vcPort(  )
       //.io_outBody_flitID(  )
       //.io_outBody_payload(  )
  );
  CreditGen CreditGen_4(
       .io_outCredit_grant( CreditGen_4_io_outCredit_grant ),
       .io_inGrant( T1134 )
  );
  RouterRegFile RouterRegFile_4(.clk(clk), .reset(reset),
       .io_writeData( T1132 ),
       .io_writeEnable( T1129 ),
       //.io_full(  )
       .io_readData( RouterRegFile_4_io_readData ),
       .io_readValid( RouterRegFile_4_io_readValid ),
       .io_readIncrement( T1116 ),
       .io_writePipelineReg_2( RouterRegFile_4_io_readPipelineReg_1 ),
       .io_writePipelineReg_1( RouterRegFile_4_io_readPipelineReg_0 ),
       .io_writePipelineReg_0( T3153 ),
       .io_wePipelineReg_2( T1105 ),
       .io_wePipelineReg_1( T1102 ),
       .io_wePipelineReg_0( T1100 ),
       //.io_readPipelineReg_2(  )
       .io_readPipelineReg_1( RouterRegFile_4_io_readPipelineReg_1 ),
       .io_readPipelineReg_0( RouterRegFile_4_io_readPipelineReg_0 ),
       //.io_rvPipelineReg_2(  )
       .io_rvPipelineReg_1( RouterRegFile_4_io_rvPipelineReg_1 ),
       .io_rvPipelineReg_0( RouterRegFile_4_io_rvPipelineReg_0 )
  );
  RouterBuffer RouterBuffer_4(.clk(clk), .reset(reset),
       .io_enq_ready( RouterBuffer_4_io_enq_ready ),
       .io_enq_valid( T1099 ),
       .io_enq_bits_x( io_inChannels_2_flit_x ),
       .io_deq_ready( T1080 ),
       .io_deq_valid( RouterBuffer_4_io_deq_valid ),
       .io_deq_bits_x( RouterBuffer_4_io_deq_bits_x )
  );
  CMeshDOR_0 CMeshDOR_4(
       .io_inHeadFlit_packetID( T1079 ),
       .io_inHeadFlit_isTail( T1078 ),
       .io_inHeadFlit_vcPort( T1077 ),
       .io_inHeadFlit_packetType( T1076 ),
       .io_inHeadFlit_destination_2( T1075 ),
       .io_inHeadFlit_destination_1( T1074 ),
       .io_inHeadFlit_destination_0( T1073 ),
       .io_inHeadFlit_priorityLevel( T1070 ),
       .io_outHeadFlit_packetID( CMeshDOR_4_io_outHeadFlit_packetID ),
       .io_outHeadFlit_isTail( CMeshDOR_4_io_outHeadFlit_isTail ),
       .io_outHeadFlit_vcPort( CMeshDOR_4_io_outHeadFlit_vcPort ),
       .io_outHeadFlit_packetType( CMeshDOR_4_io_outHeadFlit_packetType ),
       .io_outHeadFlit_destination_2( CMeshDOR_4_io_outHeadFlit_destination_2 ),
       .io_outHeadFlit_destination_1( CMeshDOR_4_io_outHeadFlit_destination_1 ),
       .io_outHeadFlit_destination_0( CMeshDOR_4_io_outHeadFlit_destination_0 ),
       .io_outHeadFlit_priorityLevel( CMeshDOR_4_io_outHeadFlit_priorityLevel ),
       .io_result( CMeshDOR_4_io_result ),
       .io_vcsAvailable_4( CMeshDOR_4_io_vcsAvailable_4 ),
       .io_vcsAvailable_3( CMeshDOR_4_io_vcsAvailable_3 ),
       .io_vcsAvailable_2( CMeshDOR_4_io_vcsAvailable_2 ),
       .io_vcsAvailable_1( CMeshDOR_4_io_vcsAvailable_1 ),
       .io_vcsAvailable_0( CMeshDOR_4_io_vcsAvailable_0 )
  );
  VCRouterStateManagement VCRouterStateManagement_4(.clk(clk), .reset(reset),
       .io_inputBufferValid( RouterBuffer_4_io_deq_valid ),
       .io_routingComplete( R1069 ),
       .io_inputBufferIsTail( T1060 ),
       .io_vcAllocGranted( vcAllocator_io_resources_4_valid ),
       .io_swAllocGranted( T1040 ),
       .io_creditsAvail( T1021 ),
       .io_outputReady( T1008 ),
       .io_currentState( VCRouterStateManagement_4_io_currentState )
  );
  ReplaceVCPort ReplaceVCPort_4(
       .io_oldFlit_x( T1006 ),
       .io_newVCPort( T3147 ),
       .io_newFlit_x( ReplaceVCPort_4_io_newFlit_x )
  );
  Flit2FlitBundle Flit2FlitBundle_4(
       .io_inFlit_x( T1000 )
       //.io_outHead_packetID(  )
       //.io_outHead_isTail(  )
       //.io_outHead_vcPort(  )
       //.io_outHead_packetType(  )
       //.io_outHead_destination_2(  )
       //.io_outHead_destination_1(  )
       //.io_outHead_destination_0(  )
       //.io_outHead_priorityLevel(  )
       //.io_outBody_packetID(  )
       //.io_outBody_isTail(  )
       //.io_outBody_vcPort(  )
       //.io_outBody_flitID(  )
       //.io_outBody_payload(  )
  );
  CreditGen CreditGen_5(
       .io_outCredit_grant( CreditGen_5_io_outCredit_grant ),
       .io_inGrant( T990 )
  );
  RouterRegFile RouterRegFile_5(.clk(clk), .reset(reset),
       .io_writeData( T988 ),
       .io_writeEnable( T985 ),
       //.io_full(  )
       .io_readData( RouterRegFile_5_io_readData ),
       .io_readValid( RouterRegFile_5_io_readValid ),
       .io_readIncrement( T972 ),
       .io_writePipelineReg_2( RouterRegFile_5_io_readPipelineReg_1 ),
       .io_writePipelineReg_1( RouterRegFile_5_io_readPipelineReg_0 ),
       .io_writePipelineReg_0( T3146 ),
       .io_wePipelineReg_2( T961 ),
       .io_wePipelineReg_1( T958 ),
       .io_wePipelineReg_0( T956 ),
       //.io_readPipelineReg_2(  )
       .io_readPipelineReg_1( RouterRegFile_5_io_readPipelineReg_1 ),
       .io_readPipelineReg_0( RouterRegFile_5_io_readPipelineReg_0 ),
       //.io_rvPipelineReg_2(  )
       .io_rvPipelineReg_1( RouterRegFile_5_io_rvPipelineReg_1 ),
       .io_rvPipelineReg_0( RouterRegFile_5_io_rvPipelineReg_0 )
  );
  RouterBuffer RouterBuffer_5(.clk(clk), .reset(reset),
       .io_enq_ready( RouterBuffer_5_io_enq_ready ),
       .io_enq_valid( T955 ),
       .io_enq_bits_x( io_inChannels_2_flit_x ),
       .io_deq_ready( T936 ),
       .io_deq_valid( RouterBuffer_5_io_deq_valid ),
       .io_deq_bits_x( RouterBuffer_5_io_deq_bits_x )
  );
  CMeshDOR_0 CMeshDOR_5(
       .io_inHeadFlit_packetID( T935 ),
       .io_inHeadFlit_isTail( T934 ),
       .io_inHeadFlit_vcPort( T933 ),
       .io_inHeadFlit_packetType( T932 ),
       .io_inHeadFlit_destination_2( T931 ),
       .io_inHeadFlit_destination_1( T930 ),
       .io_inHeadFlit_destination_0( T929 ),
       .io_inHeadFlit_priorityLevel( T926 ),
       .io_outHeadFlit_packetID( CMeshDOR_5_io_outHeadFlit_packetID ),
       .io_outHeadFlit_isTail( CMeshDOR_5_io_outHeadFlit_isTail ),
       .io_outHeadFlit_vcPort( CMeshDOR_5_io_outHeadFlit_vcPort ),
       .io_outHeadFlit_packetType( CMeshDOR_5_io_outHeadFlit_packetType ),
       .io_outHeadFlit_destination_2( CMeshDOR_5_io_outHeadFlit_destination_2 ),
       .io_outHeadFlit_destination_1( CMeshDOR_5_io_outHeadFlit_destination_1 ),
       .io_outHeadFlit_destination_0( CMeshDOR_5_io_outHeadFlit_destination_0 ),
       .io_outHeadFlit_priorityLevel( CMeshDOR_5_io_outHeadFlit_priorityLevel ),
       .io_result( CMeshDOR_5_io_result ),
       .io_vcsAvailable_4( CMeshDOR_5_io_vcsAvailable_4 ),
       .io_vcsAvailable_3( CMeshDOR_5_io_vcsAvailable_3 ),
       .io_vcsAvailable_2( CMeshDOR_5_io_vcsAvailable_2 ),
       .io_vcsAvailable_1( CMeshDOR_5_io_vcsAvailable_1 ),
       .io_vcsAvailable_0( CMeshDOR_5_io_vcsAvailable_0 )
  );
  VCRouterStateManagement VCRouterStateManagement_5(.clk(clk), .reset(reset),
       .io_inputBufferValid( RouterBuffer_5_io_deq_valid ),
       .io_routingComplete( R925 ),
       .io_inputBufferIsTail( T916 ),
       .io_vcAllocGranted( vcAllocator_io_resources_5_valid ),
       .io_swAllocGranted( T896 ),
       .io_creditsAvail( T877 ),
       .io_outputReady( T864 ),
       .io_currentState( VCRouterStateManagement_5_io_currentState )
  );
  ReplaceVCPort ReplaceVCPort_5(
       .io_oldFlit_x( T862 ),
       .io_newVCPort( T3140 ),
       .io_newFlit_x( ReplaceVCPort_5_io_newFlit_x )
  );
  Flit2FlitBundle Flit2FlitBundle_5(
       .io_inFlit_x( T856 )
       //.io_outHead_packetID(  )
       //.io_outHead_isTail(  )
       //.io_outHead_vcPort(  )
       //.io_outHead_packetType(  )
       //.io_outHead_destination_2(  )
       //.io_outHead_destination_1(  )
       //.io_outHead_destination_0(  )
       //.io_outHead_priorityLevel(  )
       //.io_outBody_packetID(  )
       //.io_outBody_isTail(  )
       //.io_outBody_vcPort(  )
       //.io_outBody_flitID(  )
       //.io_outBody_payload(  )
  );
  CreditGen CreditGen_6(
       .io_outCredit_grant( CreditGen_6_io_outCredit_grant ),
       .io_inGrant( T846 )
  );
  RouterRegFile RouterRegFile_6(.clk(clk), .reset(reset),
       .io_writeData( T844 ),
       .io_writeEnable( T841 ),
       //.io_full(  )
       .io_readData( RouterRegFile_6_io_readData ),
       .io_readValid( RouterRegFile_6_io_readValid ),
       .io_readIncrement( T828 ),
       .io_writePipelineReg_2( RouterRegFile_6_io_readPipelineReg_1 ),
       .io_writePipelineReg_1( RouterRegFile_6_io_readPipelineReg_0 ),
       .io_writePipelineReg_0( T3139 ),
       .io_wePipelineReg_2( T817 ),
       .io_wePipelineReg_1( T814 ),
       .io_wePipelineReg_0( T812 ),
       //.io_readPipelineReg_2(  )
       .io_readPipelineReg_1( RouterRegFile_6_io_readPipelineReg_1 ),
       .io_readPipelineReg_0( RouterRegFile_6_io_readPipelineReg_0 ),
       //.io_rvPipelineReg_2(  )
       .io_rvPipelineReg_1( RouterRegFile_6_io_rvPipelineReg_1 ),
       .io_rvPipelineReg_0( RouterRegFile_6_io_rvPipelineReg_0 )
  );
  RouterBuffer RouterBuffer_6(.clk(clk), .reset(reset),
       .io_enq_ready( RouterBuffer_6_io_enq_ready ),
       .io_enq_valid( T811 ),
       .io_enq_bits_x( io_inChannels_3_flit_x ),
       .io_deq_ready( T792 ),
       .io_deq_valid( RouterBuffer_6_io_deq_valid ),
       .io_deq_bits_x( RouterBuffer_6_io_deq_bits_x )
  );
  CMeshDOR_0 CMeshDOR_6(
       .io_inHeadFlit_packetID( T791 ),
       .io_inHeadFlit_isTail( T790 ),
       .io_inHeadFlit_vcPort( T789 ),
       .io_inHeadFlit_packetType( T788 ),
       .io_inHeadFlit_destination_2( T787 ),
       .io_inHeadFlit_destination_1( T786 ),
       .io_inHeadFlit_destination_0( T785 ),
       .io_inHeadFlit_priorityLevel( T782 ),
       .io_outHeadFlit_packetID( CMeshDOR_6_io_outHeadFlit_packetID ),
       .io_outHeadFlit_isTail( CMeshDOR_6_io_outHeadFlit_isTail ),
       .io_outHeadFlit_vcPort( CMeshDOR_6_io_outHeadFlit_vcPort ),
       .io_outHeadFlit_packetType( CMeshDOR_6_io_outHeadFlit_packetType ),
       .io_outHeadFlit_destination_2( CMeshDOR_6_io_outHeadFlit_destination_2 ),
       .io_outHeadFlit_destination_1( CMeshDOR_6_io_outHeadFlit_destination_1 ),
       .io_outHeadFlit_destination_0( CMeshDOR_6_io_outHeadFlit_destination_0 ),
       .io_outHeadFlit_priorityLevel( CMeshDOR_6_io_outHeadFlit_priorityLevel ),
       .io_result( CMeshDOR_6_io_result ),
       .io_vcsAvailable_4( CMeshDOR_6_io_vcsAvailable_4 ),
       .io_vcsAvailable_3( CMeshDOR_6_io_vcsAvailable_3 ),
       .io_vcsAvailable_2( CMeshDOR_6_io_vcsAvailable_2 ),
       .io_vcsAvailable_1( CMeshDOR_6_io_vcsAvailable_1 ),
       .io_vcsAvailable_0( CMeshDOR_6_io_vcsAvailable_0 )
  );
  VCRouterStateManagement VCRouterStateManagement_6(.clk(clk), .reset(reset),
       .io_inputBufferValid( RouterBuffer_6_io_deq_valid ),
       .io_routingComplete( R781 ),
       .io_inputBufferIsTail( T772 ),
       .io_vcAllocGranted( vcAllocator_io_resources_6_valid ),
       .io_swAllocGranted( T752 ),
       .io_creditsAvail( T733 ),
       .io_outputReady( T720 ),
       .io_currentState( VCRouterStateManagement_6_io_currentState )
  );
  ReplaceVCPort ReplaceVCPort_6(
       .io_oldFlit_x( T718 ),
       .io_newVCPort( T3133 ),
       .io_newFlit_x( ReplaceVCPort_6_io_newFlit_x )
  );
  Flit2FlitBundle Flit2FlitBundle_6(
       .io_inFlit_x( T712 )
       //.io_outHead_packetID(  )
       //.io_outHead_isTail(  )
       //.io_outHead_vcPort(  )
       //.io_outHead_packetType(  )
       //.io_outHead_destination_2(  )
       //.io_outHead_destination_1(  )
       //.io_outHead_destination_0(  )
       //.io_outHead_priorityLevel(  )
       //.io_outBody_packetID(  )
       //.io_outBody_isTail(  )
       //.io_outBody_vcPort(  )
       //.io_outBody_flitID(  )
       //.io_outBody_payload(  )
  );
  CreditGen CreditGen_7(
       .io_outCredit_grant( CreditGen_7_io_outCredit_grant ),
       .io_inGrant( T702 )
  );
  RouterRegFile RouterRegFile_7(.clk(clk), .reset(reset),
       .io_writeData( T700 ),
       .io_writeEnable( T697 ),
       //.io_full(  )
       .io_readData( RouterRegFile_7_io_readData ),
       .io_readValid( RouterRegFile_7_io_readValid ),
       .io_readIncrement( T684 ),
       .io_writePipelineReg_2( RouterRegFile_7_io_readPipelineReg_1 ),
       .io_writePipelineReg_1( RouterRegFile_7_io_readPipelineReg_0 ),
       .io_writePipelineReg_0( T3132 ),
       .io_wePipelineReg_2( T673 ),
       .io_wePipelineReg_1( T670 ),
       .io_wePipelineReg_0( T668 ),
       //.io_readPipelineReg_2(  )
       .io_readPipelineReg_1( RouterRegFile_7_io_readPipelineReg_1 ),
       .io_readPipelineReg_0( RouterRegFile_7_io_readPipelineReg_0 ),
       //.io_rvPipelineReg_2(  )
       .io_rvPipelineReg_1( RouterRegFile_7_io_rvPipelineReg_1 ),
       .io_rvPipelineReg_0( RouterRegFile_7_io_rvPipelineReg_0 )
  );
  RouterBuffer RouterBuffer_7(.clk(clk), .reset(reset),
       .io_enq_ready( RouterBuffer_7_io_enq_ready ),
       .io_enq_valid( T667 ),
       .io_enq_bits_x( io_inChannels_3_flit_x ),
       .io_deq_ready( T648 ),
       .io_deq_valid( RouterBuffer_7_io_deq_valid ),
       .io_deq_bits_x( RouterBuffer_7_io_deq_bits_x )
  );
  CMeshDOR_0 CMeshDOR_7(
       .io_inHeadFlit_packetID( T647 ),
       .io_inHeadFlit_isTail( T646 ),
       .io_inHeadFlit_vcPort( T645 ),
       .io_inHeadFlit_packetType( T644 ),
       .io_inHeadFlit_destination_2( T643 ),
       .io_inHeadFlit_destination_1( T642 ),
       .io_inHeadFlit_destination_0( T641 ),
       .io_inHeadFlit_priorityLevel( T638 ),
       .io_outHeadFlit_packetID( CMeshDOR_7_io_outHeadFlit_packetID ),
       .io_outHeadFlit_isTail( CMeshDOR_7_io_outHeadFlit_isTail ),
       .io_outHeadFlit_vcPort( CMeshDOR_7_io_outHeadFlit_vcPort ),
       .io_outHeadFlit_packetType( CMeshDOR_7_io_outHeadFlit_packetType ),
       .io_outHeadFlit_destination_2( CMeshDOR_7_io_outHeadFlit_destination_2 ),
       .io_outHeadFlit_destination_1( CMeshDOR_7_io_outHeadFlit_destination_1 ),
       .io_outHeadFlit_destination_0( CMeshDOR_7_io_outHeadFlit_destination_0 ),
       .io_outHeadFlit_priorityLevel( CMeshDOR_7_io_outHeadFlit_priorityLevel ),
       .io_result( CMeshDOR_7_io_result ),
       .io_vcsAvailable_4( CMeshDOR_7_io_vcsAvailable_4 ),
       .io_vcsAvailable_3( CMeshDOR_7_io_vcsAvailable_3 ),
       .io_vcsAvailable_2( CMeshDOR_7_io_vcsAvailable_2 ),
       .io_vcsAvailable_1( CMeshDOR_7_io_vcsAvailable_1 ),
       .io_vcsAvailable_0( CMeshDOR_7_io_vcsAvailable_0 )
  );
  VCRouterStateManagement VCRouterStateManagement_7(.clk(clk), .reset(reset),
       .io_inputBufferValid( RouterBuffer_7_io_deq_valid ),
       .io_routingComplete( R637 ),
       .io_inputBufferIsTail( T628 ),
       .io_vcAllocGranted( vcAllocator_io_resources_7_valid ),
       .io_swAllocGranted( T608 ),
       .io_creditsAvail( T589 ),
       .io_outputReady( T576 ),
       .io_currentState( VCRouterStateManagement_7_io_currentState )
  );
  ReplaceVCPort ReplaceVCPort_7(
       .io_oldFlit_x( T574 ),
       .io_newVCPort( T3126 ),
       .io_newFlit_x( ReplaceVCPort_7_io_newFlit_x )
  );
  Flit2FlitBundle Flit2FlitBundle_7(
       .io_inFlit_x( T568 )
       //.io_outHead_packetID(  )
       //.io_outHead_isTail(  )
       //.io_outHead_vcPort(  )
       //.io_outHead_packetType(  )
       //.io_outHead_destination_2(  )
       //.io_outHead_destination_1(  )
       //.io_outHead_destination_0(  )
       //.io_outHead_priorityLevel(  )
       //.io_outBody_packetID(  )
       //.io_outBody_isTail(  )
       //.io_outBody_vcPort(  )
       //.io_outBody_flitID(  )
       //.io_outBody_payload(  )
  );
  CreditGen CreditGen_8(
       .io_outCredit_grant( CreditGen_8_io_outCredit_grant ),
       .io_inGrant( T558 )
  );
  RouterRegFile RouterRegFile_8(.clk(clk), .reset(reset),
       .io_writeData( T556 ),
       .io_writeEnable( T553 ),
       //.io_full(  )
       .io_readData( RouterRegFile_8_io_readData ),
       .io_readValid( RouterRegFile_8_io_readValid ),
       .io_readIncrement( T540 ),
       .io_writePipelineReg_2( RouterRegFile_8_io_readPipelineReg_1 ),
       .io_writePipelineReg_1( RouterRegFile_8_io_readPipelineReg_0 ),
       .io_writePipelineReg_0( T3125 ),
       .io_wePipelineReg_2( T529 ),
       .io_wePipelineReg_1( T526 ),
       .io_wePipelineReg_0( T524 ),
       //.io_readPipelineReg_2(  )
       .io_readPipelineReg_1( RouterRegFile_8_io_readPipelineReg_1 ),
       .io_readPipelineReg_0( RouterRegFile_8_io_readPipelineReg_0 ),
       //.io_rvPipelineReg_2(  )
       .io_rvPipelineReg_1( RouterRegFile_8_io_rvPipelineReg_1 ),
       .io_rvPipelineReg_0( RouterRegFile_8_io_rvPipelineReg_0 )
  );
  RouterBuffer RouterBuffer_8(.clk(clk), .reset(reset),
       .io_enq_ready( RouterBuffer_8_io_enq_ready ),
       .io_enq_valid( T523 ),
       .io_enq_bits_x( io_inChannels_4_flit_x ),
       .io_deq_ready( T504 ),
       .io_deq_valid( RouterBuffer_8_io_deq_valid ),
       .io_deq_bits_x( RouterBuffer_8_io_deq_bits_x )
  );
  CMeshDOR_0 CMeshDOR_8(
       .io_inHeadFlit_packetID( T503 ),
       .io_inHeadFlit_isTail( T502 ),
       .io_inHeadFlit_vcPort( T501 ),
       .io_inHeadFlit_packetType( T500 ),
       .io_inHeadFlit_destination_2( T499 ),
       .io_inHeadFlit_destination_1( T498 ),
       .io_inHeadFlit_destination_0( T497 ),
       .io_inHeadFlit_priorityLevel( T494 ),
       .io_outHeadFlit_packetID( CMeshDOR_8_io_outHeadFlit_packetID ),
       .io_outHeadFlit_isTail( CMeshDOR_8_io_outHeadFlit_isTail ),
       .io_outHeadFlit_vcPort( CMeshDOR_8_io_outHeadFlit_vcPort ),
       .io_outHeadFlit_packetType( CMeshDOR_8_io_outHeadFlit_packetType ),
       .io_outHeadFlit_destination_2( CMeshDOR_8_io_outHeadFlit_destination_2 ),
       .io_outHeadFlit_destination_1( CMeshDOR_8_io_outHeadFlit_destination_1 ),
       .io_outHeadFlit_destination_0( CMeshDOR_8_io_outHeadFlit_destination_0 ),
       .io_outHeadFlit_priorityLevel( CMeshDOR_8_io_outHeadFlit_priorityLevel ),
       .io_result( CMeshDOR_8_io_result ),
       .io_vcsAvailable_4( CMeshDOR_8_io_vcsAvailable_4 ),
       .io_vcsAvailable_3( CMeshDOR_8_io_vcsAvailable_3 ),
       .io_vcsAvailable_2( CMeshDOR_8_io_vcsAvailable_2 ),
       .io_vcsAvailable_1( CMeshDOR_8_io_vcsAvailable_1 ),
       .io_vcsAvailable_0( CMeshDOR_8_io_vcsAvailable_0 )
  );
  VCRouterStateManagement VCRouterStateManagement_8(.clk(clk), .reset(reset),
       .io_inputBufferValid( RouterBuffer_8_io_deq_valid ),
       .io_routingComplete( R493 ),
       .io_inputBufferIsTail( T484 ),
       .io_vcAllocGranted( vcAllocator_io_resources_8_valid ),
       .io_swAllocGranted( T464 ),
       .io_creditsAvail( T445 ),
       .io_outputReady( T432 ),
       .io_currentState( VCRouterStateManagement_8_io_currentState )
  );
  ReplaceVCPort ReplaceVCPort_8(
       .io_oldFlit_x( T430 ),
       .io_newVCPort( T3119 ),
       .io_newFlit_x( ReplaceVCPort_8_io_newFlit_x )
  );
  Flit2FlitBundle Flit2FlitBundle_8(
       .io_inFlit_x( T424 )
       //.io_outHead_packetID(  )
       //.io_outHead_isTail(  )
       //.io_outHead_vcPort(  )
       //.io_outHead_packetType(  )
       //.io_outHead_destination_2(  )
       //.io_outHead_destination_1(  )
       //.io_outHead_destination_0(  )
       //.io_outHead_priorityLevel(  )
       //.io_outBody_packetID(  )
       //.io_outBody_isTail(  )
       //.io_outBody_vcPort(  )
       //.io_outBody_flitID(  )
       //.io_outBody_payload(  )
  );
  CreditGen CreditGen_9(
       .io_outCredit_grant( CreditGen_9_io_outCredit_grant ),
       .io_inGrant( T414 )
  );
  RouterRegFile RouterRegFile_9(.clk(clk), .reset(reset),
       .io_writeData( T412 ),
       .io_writeEnable( T409 ),
       //.io_full(  )
       .io_readData( RouterRegFile_9_io_readData ),
       .io_readValid( RouterRegFile_9_io_readValid ),
       .io_readIncrement( T396 ),
       .io_writePipelineReg_2( RouterRegFile_9_io_readPipelineReg_1 ),
       .io_writePipelineReg_1( RouterRegFile_9_io_readPipelineReg_0 ),
       .io_writePipelineReg_0( T3118 ),
       .io_wePipelineReg_2( T385 ),
       .io_wePipelineReg_1( T382 ),
       .io_wePipelineReg_0( T380 ),
       //.io_readPipelineReg_2(  )
       .io_readPipelineReg_1( RouterRegFile_9_io_readPipelineReg_1 ),
       .io_readPipelineReg_0( RouterRegFile_9_io_readPipelineReg_0 ),
       //.io_rvPipelineReg_2(  )
       .io_rvPipelineReg_1( RouterRegFile_9_io_rvPipelineReg_1 ),
       .io_rvPipelineReg_0( RouterRegFile_9_io_rvPipelineReg_0 )
  );
  RouterBuffer RouterBuffer_9(.clk(clk), .reset(reset),
       .io_enq_ready( RouterBuffer_9_io_enq_ready ),
       .io_enq_valid( T379 ),
       .io_enq_bits_x( io_inChannels_4_flit_x ),
       .io_deq_ready( T360 ),
       .io_deq_valid( RouterBuffer_9_io_deq_valid ),
       .io_deq_bits_x( RouterBuffer_9_io_deq_bits_x )
  );
  CMeshDOR_0 CMeshDOR_9(
       .io_inHeadFlit_packetID( T359 ),
       .io_inHeadFlit_isTail( T358 ),
       .io_inHeadFlit_vcPort( T357 ),
       .io_inHeadFlit_packetType( T356 ),
       .io_inHeadFlit_destination_2( T355 ),
       .io_inHeadFlit_destination_1( T354 ),
       .io_inHeadFlit_destination_0( T353 ),
       .io_inHeadFlit_priorityLevel( T350 ),
       .io_outHeadFlit_packetID( CMeshDOR_9_io_outHeadFlit_packetID ),
       .io_outHeadFlit_isTail( CMeshDOR_9_io_outHeadFlit_isTail ),
       .io_outHeadFlit_vcPort( CMeshDOR_9_io_outHeadFlit_vcPort ),
       .io_outHeadFlit_packetType( CMeshDOR_9_io_outHeadFlit_packetType ),
       .io_outHeadFlit_destination_2( CMeshDOR_9_io_outHeadFlit_destination_2 ),
       .io_outHeadFlit_destination_1( CMeshDOR_9_io_outHeadFlit_destination_1 ),
       .io_outHeadFlit_destination_0( CMeshDOR_9_io_outHeadFlit_destination_0 ),
       .io_outHeadFlit_priorityLevel( CMeshDOR_9_io_outHeadFlit_priorityLevel ),
       .io_result( CMeshDOR_9_io_result ),
       .io_vcsAvailable_4( CMeshDOR_9_io_vcsAvailable_4 ),
       .io_vcsAvailable_3( CMeshDOR_9_io_vcsAvailable_3 ),
       .io_vcsAvailable_2( CMeshDOR_9_io_vcsAvailable_2 ),
       .io_vcsAvailable_1( CMeshDOR_9_io_vcsAvailable_1 ),
       .io_vcsAvailable_0( CMeshDOR_9_io_vcsAvailable_0 )
  );
  VCRouterStateManagement VCRouterStateManagement_9(.clk(clk), .reset(reset),
       .io_inputBufferValid( RouterBuffer_9_io_deq_valid ),
       .io_routingComplete( R349 ),
       .io_inputBufferIsTail( T340 ),
       .io_vcAllocGranted( vcAllocator_io_resources_9_valid ),
       .io_swAllocGranted( T320 ),
       .io_creditsAvail( T301 ),
       .io_outputReady( T288 ),
       .io_currentState( VCRouterStateManagement_9_io_currentState )
  );
  ReplaceVCPort ReplaceVCPort_9(
       .io_oldFlit_x( T286 ),
       .io_newVCPort( T3112 ),
       .io_newFlit_x( ReplaceVCPort_9_io_newFlit_x )
  );
  Flit2FlitBundle Flit2FlitBundle_9(
       .io_inFlit_x( T280 )
       //.io_outHead_packetID(  )
       //.io_outHead_isTail(  )
       //.io_outHead_vcPort(  )
       //.io_outHead_packetType(  )
       //.io_outHead_destination_2(  )
       //.io_outHead_destination_1(  )
       //.io_outHead_destination_0(  )
       //.io_outHead_priorityLevel(  )
       //.io_outBody_packetID(  )
       //.io_outBody_isTail(  )
       //.io_outBody_vcPort(  )
       //.io_outBody_flitID(  )
       //.io_outBody_payload(  )
  );
  CreditCon CreditCon(.clk(clk), .reset(reset),
       .io_inCredit_grant( io_outChannels_0_credit_0_grant ),
       .io_inConsume( T278 ),
       .io_outCredit( CreditCon_io_outCredit )
       //.io_almostOut(  )
  );
  CreditCon CreditCon_1(.clk(clk), .reset(reset),
       .io_inCredit_grant( io_outChannels_0_credit_1_grant ),
       .io_inConsume( T268 ),
       .io_outCredit( CreditCon_1_io_outCredit )
       //.io_almostOut(  )
  );
  MuxN_1 MuxN(
       //.io_ins_1(  )
       //.io_ins_0(  )
       //.io_sel(  )
       //.io_out(  )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign MuxN.io_ins_1 = {1{1'b0}};
    assign MuxN.io_ins_0 = {1{1'b0}};
    assign MuxN.io_sel = {1{1'b0}};
// synthesis translate_on
`endif
  CreditCon CreditCon_2(.clk(clk), .reset(reset),
       .io_inCredit_grant( io_outChannels_1_credit_0_grant ),
       .io_inConsume( T266 ),
       .io_outCredit( CreditCon_2_io_outCredit )
       //.io_almostOut(  )
  );
  CreditCon CreditCon_3(.clk(clk), .reset(reset),
       .io_inCredit_grant( io_outChannels_1_credit_1_grant ),
       .io_inConsume( T256 ),
       .io_outCredit( CreditCon_3_io_outCredit )
       //.io_almostOut(  )
  );
  MuxN_1 MuxN_1(
       //.io_ins_1(  )
       //.io_ins_0(  )
       //.io_sel(  )
       //.io_out(  )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign MuxN_1.io_ins_1 = {1{1'b0}};
    assign MuxN_1.io_ins_0 = {1{1'b0}};
    assign MuxN_1.io_sel = {1{1'b0}};
// synthesis translate_on
`endif
  CreditCon CreditCon_4(.clk(clk), .reset(reset),
       .io_inCredit_grant( io_outChannels_2_credit_0_grant ),
       .io_inConsume( T254 ),
       .io_outCredit( CreditCon_4_io_outCredit )
       //.io_almostOut(  )
  );
  CreditCon CreditCon_5(.clk(clk), .reset(reset),
       .io_inCredit_grant( io_outChannels_2_credit_1_grant ),
       .io_inConsume( T244 ),
       .io_outCredit( CreditCon_5_io_outCredit )
       //.io_almostOut(  )
  );
  MuxN_1 MuxN_2(
       //.io_ins_1(  )
       //.io_ins_0(  )
       //.io_sel(  )
       //.io_out(  )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign MuxN_2.io_ins_1 = {1{1'b0}};
    assign MuxN_2.io_ins_0 = {1{1'b0}};
    assign MuxN_2.io_sel = {1{1'b0}};
// synthesis translate_on
`endif
  CreditCon CreditCon_6(.clk(clk), .reset(reset),
       .io_inCredit_grant( io_outChannels_3_credit_0_grant ),
       .io_inConsume( T242 ),
       .io_outCredit( CreditCon_6_io_outCredit )
       //.io_almostOut(  )
  );
  CreditCon CreditCon_7(.clk(clk), .reset(reset),
       .io_inCredit_grant( io_outChannels_3_credit_1_grant ),
       .io_inConsume( T232 ),
       .io_outCredit( CreditCon_7_io_outCredit )
       //.io_almostOut(  )
  );
  MuxN_1 MuxN_3(
       //.io_ins_1(  )
       //.io_ins_0(  )
       //.io_sel(  )
       //.io_out(  )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign MuxN_3.io_ins_1 = {1{1'b0}};
    assign MuxN_3.io_ins_0 = {1{1'b0}};
    assign MuxN_3.io_sel = {1{1'b0}};
// synthesis translate_on
`endif
  CreditCon CreditCon_8(.clk(clk), .reset(reset),
       .io_inCredit_grant( io_outChannels_4_credit_0_grant ),
       .io_inConsume( T230 ),
       .io_outCredit( CreditCon_8_io_outCredit )
       //.io_almostOut(  )
  );
  CreditCon CreditCon_9(.clk(clk), .reset(reset),
       .io_inCredit_grant( io_outChannels_4_credit_1_grant ),
       .io_inConsume( T220 ),
       .io_outCredit( CreditCon_9_io_outCredit )
       //.io_almostOut(  )
  );
  MuxN_1 MuxN_4(
       //.io_ins_1(  )
       //.io_ins_0(  )
       //.io_sel(  )
       //.io_out(  )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign MuxN_4.io_ins_1 = {1{1'b0}};
    assign MuxN_4.io_ins_0 = {1{1'b0}};
    assign MuxN_4.io_sel = {1{1'b0}};
// synthesis translate_on
`endif

  always @(posedge clk) begin
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T215 <= 1'b1;
  if(!T216 && T215 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "SimpleVCRouter: Flit with VC port/*? in < (class OpenSoC.SimpleVCRouter)>*/ Chisel.UInt(width=1, connect to 1 inputs: ([Chisel.Mux] in OpenSoC.SimpleVCRouter)) attempting to write to VC 0");
    $finish;
  end
// synthesis translate_on
`endif
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T198 <= 1'b1;
  if(!T199 && T198 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "SimpleVCRouter:Vector(0, 0) Insufficent space in input buffer - Credit Ready asserted when Routing In Buffer not ready inputPort= 0 curVC = 0");
    $finish;
  end
// synthesis translate_on
`endif
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T193 <= 1'b1;
  if(!T194 && T193 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "SimpleVCRouter: Flit with VC port/*? in < (class OpenSoC.SimpleVCRouter)>*/ Chisel.UInt(width=1, connect to 1 inputs: ([Chisel.Mux] in OpenSoC.SimpleVCRouter)) attempting to write to VC 1");
    $finish;
  end
// synthesis translate_on
`endif
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T176 <= 1'b1;
  if(!T177 && T176 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "SimpleVCRouter:Vector(0, 0) Insufficent space in input buffer - Credit Ready asserted when Routing In Buffer not ready inputPort= 0 curVC = 1");
    $finish;
  end
// synthesis translate_on
`endif
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T171 <= 1'b1;
  if(!T172 && T171 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "SimpleVCRouter: Flit with VC port/*? in < (class OpenSoC.SimpleVCRouter)>*/ Chisel.UInt(width=1, connect to 1 inputs: ([Chisel.Mux] in OpenSoC.SimpleVCRouter)) attempting to write to VC 0");
    $finish;
  end
// synthesis translate_on
`endif
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T154 <= 1'b1;
  if(!T155 && T154 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "SimpleVCRouter:Vector(0, 0) Insufficent space in input buffer - Credit Ready asserted when Routing In Buffer not ready inputPort= 1 curVC = 0");
    $finish;
  end
// synthesis translate_on
`endif
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T149 <= 1'b1;
  if(!T150 && T149 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "SimpleVCRouter: Flit with VC port/*? in < (class OpenSoC.SimpleVCRouter)>*/ Chisel.UInt(width=1, connect to 1 inputs: ([Chisel.Mux] in OpenSoC.SimpleVCRouter)) attempting to write to VC 1");
    $finish;
  end
// synthesis translate_on
`endif
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T132 <= 1'b1;
  if(!T133 && T132 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "SimpleVCRouter:Vector(0, 0) Insufficent space in input buffer - Credit Ready asserted when Routing In Buffer not ready inputPort= 1 curVC = 1");
    $finish;
  end
// synthesis translate_on
`endif
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T127 <= 1'b1;
  if(!T128 && T127 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "SimpleVCRouter: Flit with VC port/*? in < (class OpenSoC.SimpleVCRouter)>*/ Chisel.UInt(width=1, connect to 1 inputs: ([Chisel.Mux] in OpenSoC.SimpleVCRouter)) attempting to write to VC 0");
    $finish;
  end
// synthesis translate_on
`endif
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T110 <= 1'b1;
  if(!T111 && T110 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "SimpleVCRouter:Vector(0, 0) Insufficent space in input buffer - Credit Ready asserted when Routing In Buffer not ready inputPort= 2 curVC = 0");
    $finish;
  end
// synthesis translate_on
`endif
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T105 <= 1'b1;
  if(!T106 && T105 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "SimpleVCRouter: Flit with VC port/*? in < (class OpenSoC.SimpleVCRouter)>*/ Chisel.UInt(width=1, connect to 1 inputs: ([Chisel.Mux] in OpenSoC.SimpleVCRouter)) attempting to write to VC 1");
    $finish;
  end
// synthesis translate_on
`endif
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T88 <= 1'b1;
  if(!T89 && T88 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "SimpleVCRouter:Vector(0, 0) Insufficent space in input buffer - Credit Ready asserted when Routing In Buffer not ready inputPort= 2 curVC = 1");
    $finish;
  end
// synthesis translate_on
`endif
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T83 <= 1'b1;
  if(!T84 && T83 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "SimpleVCRouter: Flit with VC port/*? in < (class OpenSoC.SimpleVCRouter)>*/ Chisel.UInt(width=1, connect to 1 inputs: ([Chisel.Mux] in OpenSoC.SimpleVCRouter)) attempting to write to VC 0");
    $finish;
  end
// synthesis translate_on
`endif
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T66 <= 1'b1;
  if(!T67 && T66 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "SimpleVCRouter:Vector(0, 0) Insufficent space in input buffer - Credit Ready asserted when Routing In Buffer not ready inputPort= 3 curVC = 0");
    $finish;
  end
// synthesis translate_on
`endif
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T61 <= 1'b1;
  if(!T62 && T61 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "SimpleVCRouter: Flit with VC port/*? in < (class OpenSoC.SimpleVCRouter)>*/ Chisel.UInt(width=1, connect to 1 inputs: ([Chisel.Mux] in OpenSoC.SimpleVCRouter)) attempting to write to VC 1");
    $finish;
  end
// synthesis translate_on
`endif
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T44 <= 1'b1;
  if(!T45 && T44 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "SimpleVCRouter:Vector(0, 0) Insufficent space in input buffer - Credit Ready asserted when Routing In Buffer not ready inputPort= 3 curVC = 1");
    $finish;
  end
// synthesis translate_on
`endif
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T39 <= 1'b1;
  if(!T40 && T39 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "SimpleVCRouter: Flit with VC port/*? in < (class OpenSoC.SimpleVCRouter)>*/ Chisel.UInt(width=1, connect to 1 inputs: ([Chisel.Mux] in OpenSoC.SimpleVCRouter)) attempting to write to VC 0");
    $finish;
  end
// synthesis translate_on
`endif
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T22 <= 1'b1;
  if(!T23 && T22 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "SimpleVCRouter:Vector(0, 0) Insufficent space in input buffer - Credit Ready asserted when Routing In Buffer not ready inputPort= 4 curVC = 0");
    $finish;
  end
// synthesis translate_on
`endif
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T17 <= 1'b1;
  if(!T18 && T17 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "SimpleVCRouter: Flit with VC port/*? in < (class OpenSoC.SimpleVCRouter)>*/ Chisel.UInt(width=1, connect to 1 inputs: ([Chisel.Mux] in OpenSoC.SimpleVCRouter)) attempting to write to VC 1");
    $finish;
  end
// synthesis translate_on
`endif
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T0 <= 1'b1;
  if(!T1 && T0 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "SimpleVCRouter:Vector(0, 0) Insufficent space in input buffer - Credit Ready asserted when Routing In Buffer not ready inputPort= 4 curVC = 1");
    $finish;
  end
// synthesis translate_on
`endif
    if(reset) begin
      R282 <= 55'h0;
    end else if(T284) begin
      R282 <= T3114;
    end
    if(reset) begin
      R295 <= 3'h0;
    end else begin
      R295 <= CMeshDOR_9_io_result;
    end
    if(reset) begin
      R349 <= 1'h0;
    end else begin
      R349 <= RouterBuffer_9_io_deq_valid;
    end
    if(reset) begin
      R426 <= 55'h0;
    end else if(T428) begin
      R426 <= T3121;
    end
    if(reset) begin
      R439 <= 3'h0;
    end else begin
      R439 <= CMeshDOR_8_io_result;
    end
    if(reset) begin
      R493 <= 1'h0;
    end else begin
      R493 <= RouterBuffer_8_io_deq_valid;
    end
    if(reset) begin
      R570 <= 55'h0;
    end else if(T572) begin
      R570 <= T3128;
    end
    if(reset) begin
      R583 <= 3'h0;
    end else begin
      R583 <= CMeshDOR_7_io_result;
    end
    if(reset) begin
      R637 <= 1'h0;
    end else begin
      R637 <= RouterBuffer_7_io_deq_valid;
    end
    if(reset) begin
      R714 <= 55'h0;
    end else if(T716) begin
      R714 <= T3135;
    end
    if(reset) begin
      R727 <= 3'h0;
    end else begin
      R727 <= CMeshDOR_6_io_result;
    end
    if(reset) begin
      R781 <= 1'h0;
    end else begin
      R781 <= RouterBuffer_6_io_deq_valid;
    end
    if(reset) begin
      R858 <= 55'h0;
    end else if(T860) begin
      R858 <= T3142;
    end
    if(reset) begin
      R871 <= 3'h0;
    end else begin
      R871 <= CMeshDOR_5_io_result;
    end
    if(reset) begin
      R925 <= 1'h0;
    end else begin
      R925 <= RouterBuffer_5_io_deq_valid;
    end
    if(reset) begin
      R1002 <= 55'h0;
    end else if(T1004) begin
      R1002 <= T3149;
    end
    if(reset) begin
      R1015 <= 3'h0;
    end else begin
      R1015 <= CMeshDOR_4_io_result;
    end
    if(reset) begin
      R1069 <= 1'h0;
    end else begin
      R1069 <= RouterBuffer_4_io_deq_valid;
    end
    if(reset) begin
      R1146 <= 55'h0;
    end else if(T1148) begin
      R1146 <= T3156;
    end
    if(reset) begin
      R1159 <= 3'h0;
    end else begin
      R1159 <= CMeshDOR_3_io_result;
    end
    if(reset) begin
      R1213 <= 1'h0;
    end else begin
      R1213 <= RouterBuffer_3_io_deq_valid;
    end
    if(reset) begin
      R1290 <= 55'h0;
    end else if(T1292) begin
      R1290 <= T3163;
    end
    if(reset) begin
      R1303 <= 3'h0;
    end else begin
      R1303 <= CMeshDOR_2_io_result;
    end
    if(reset) begin
      R1357 <= 1'h0;
    end else begin
      R1357 <= RouterBuffer_2_io_deq_valid;
    end
    if(reset) begin
      R1434 <= 55'h0;
    end else if(T1436) begin
      R1434 <= T3170;
    end
    if(reset) begin
      R1447 <= 3'h0;
    end else begin
      R1447 <= CMeshDOR_1_io_result;
    end
    if(reset) begin
      R1501 <= 1'h0;
    end else begin
      R1501 <= RouterBuffer_1_io_deq_valid;
    end
    if(reset) begin
      R1578 <= 55'h0;
    end else if(T1580) begin
      R1578 <= T3177;
    end
    if(reset) begin
      R1591 <= 3'h0;
    end else begin
      R1591 <= CMeshDOR_io_result;
    end
    if(reset) begin
      R1645 <= 1'h0;
    end else begin
      R1645 <= RouterBuffer_io_deq_valid;
    end
    validVCs_0_0 <= CMeshDOR_io_vcsAvailable_0;
    R2176 <= T2177;
    R2181 <= T2182;
    validVCs_0_1 <= CMeshDOR_io_vcsAvailable_1;
    R2186 <= T2187;
    R2191 <= T2192;
    validVCs_0_2 <= CMeshDOR_io_vcsAvailable_2;
    R2196 <= T2197;
    R2201 <= T2202;
    validVCs_0_3 <= CMeshDOR_io_vcsAvailable_3;
    R2206 <= T2207;
    R2211 <= T2212;
    validVCs_0_4 <= CMeshDOR_io_vcsAvailable_4;
    R2216 <= T2217;
    R2221 <= T2222;
    validVCs_1_0 <= CMeshDOR_1_io_vcsAvailable_0;
    R2226 <= T2227;
    R2231 <= T2232;
    validVCs_1_1 <= CMeshDOR_1_io_vcsAvailable_1;
    R2236 <= T2237;
    R2241 <= T2242;
    validVCs_1_2 <= CMeshDOR_1_io_vcsAvailable_2;
    R2246 <= T2247;
    R2251 <= T2252;
    validVCs_1_3 <= CMeshDOR_1_io_vcsAvailable_3;
    R2256 <= T2257;
    R2261 <= T2262;
    validVCs_1_4 <= CMeshDOR_1_io_vcsAvailable_4;
    R2266 <= T2267;
    R2271 <= T2272;
    validVCs_2_0 <= CMeshDOR_2_io_vcsAvailable_0;
    R2276 <= T2277;
    R2281 <= T2282;
    validVCs_2_1 <= CMeshDOR_2_io_vcsAvailable_1;
    R2286 <= T2287;
    R2291 <= T2292;
    validVCs_2_2 <= CMeshDOR_2_io_vcsAvailable_2;
    R2296 <= T2297;
    R2301 <= T2302;
    validVCs_2_3 <= CMeshDOR_2_io_vcsAvailable_3;
    R2306 <= T2307;
    R2311 <= T2312;
    validVCs_2_4 <= CMeshDOR_2_io_vcsAvailable_4;
    R2316 <= T2317;
    R2321 <= T2322;
    validVCs_3_0 <= CMeshDOR_3_io_vcsAvailable_0;
    R2326 <= T2327;
    R2331 <= T2332;
    validVCs_3_1 <= CMeshDOR_3_io_vcsAvailable_1;
    R2336 <= T2337;
    R2341 <= T2342;
    validVCs_3_2 <= CMeshDOR_3_io_vcsAvailable_2;
    R2346 <= T2347;
    R2351 <= T2352;
    validVCs_3_3 <= CMeshDOR_3_io_vcsAvailable_3;
    R2356 <= T2357;
    R2361 <= T2362;
    validVCs_3_4 <= CMeshDOR_3_io_vcsAvailable_4;
    R2366 <= T2367;
    R2371 <= T2372;
    validVCs_4_0 <= CMeshDOR_4_io_vcsAvailable_0;
    R2376 <= T2377;
    R2381 <= T2382;
    validVCs_4_1 <= CMeshDOR_4_io_vcsAvailable_1;
    R2386 <= T2387;
    R2391 <= T2392;
    validVCs_4_2 <= CMeshDOR_4_io_vcsAvailable_2;
    R2396 <= T2397;
    R2401 <= T2402;
    validVCs_4_3 <= CMeshDOR_4_io_vcsAvailable_3;
    R2406 <= T2407;
    R2411 <= T2412;
    validVCs_4_4 <= CMeshDOR_4_io_vcsAvailable_4;
    R2416 <= T2417;
    R2421 <= T2422;
    validVCs_5_0 <= CMeshDOR_5_io_vcsAvailable_0;
    R2426 <= T2427;
    R2431 <= T2432;
    validVCs_5_1 <= CMeshDOR_5_io_vcsAvailable_1;
    R2436 <= T2437;
    R2441 <= T2442;
    validVCs_5_2 <= CMeshDOR_5_io_vcsAvailable_2;
    R2446 <= T2447;
    R2451 <= T2452;
    validVCs_5_3 <= CMeshDOR_5_io_vcsAvailable_3;
    R2456 <= T2457;
    R2461 <= T2462;
    validVCs_5_4 <= CMeshDOR_5_io_vcsAvailable_4;
    R2466 <= T2467;
    R2471 <= T2472;
    validVCs_6_0 <= CMeshDOR_6_io_vcsAvailable_0;
    R2476 <= T2477;
    R2481 <= T2482;
    validVCs_6_1 <= CMeshDOR_6_io_vcsAvailable_1;
    R2486 <= T2487;
    R2491 <= T2492;
    validVCs_6_2 <= CMeshDOR_6_io_vcsAvailable_2;
    R2496 <= T2497;
    R2501 <= T2502;
    validVCs_6_3 <= CMeshDOR_6_io_vcsAvailable_3;
    R2506 <= T2507;
    R2511 <= T2512;
    validVCs_6_4 <= CMeshDOR_6_io_vcsAvailable_4;
    R2516 <= T2517;
    R2521 <= T2522;
    validVCs_7_0 <= CMeshDOR_7_io_vcsAvailable_0;
    R2526 <= T2527;
    R2531 <= T2532;
    validVCs_7_1 <= CMeshDOR_7_io_vcsAvailable_1;
    R2536 <= T2537;
    R2541 <= T2542;
    validVCs_7_2 <= CMeshDOR_7_io_vcsAvailable_2;
    R2546 <= T2547;
    R2551 <= T2552;
    validVCs_7_3 <= CMeshDOR_7_io_vcsAvailable_3;
    R2556 <= T2557;
    R2561 <= T2562;
    validVCs_7_4 <= CMeshDOR_7_io_vcsAvailable_4;
    R2566 <= T2567;
    R2571 <= T2572;
    validVCs_8_0 <= CMeshDOR_8_io_vcsAvailable_0;
    R2576 <= T2577;
    R2581 <= T2582;
    validVCs_8_1 <= CMeshDOR_8_io_vcsAvailable_1;
    R2586 <= T2587;
    R2591 <= T2592;
    validVCs_8_2 <= CMeshDOR_8_io_vcsAvailable_2;
    R2596 <= T2597;
    R2601 <= T2602;
    validVCs_8_3 <= CMeshDOR_8_io_vcsAvailable_3;
    R2606 <= T2607;
    R2611 <= T2612;
    validVCs_8_4 <= CMeshDOR_8_io_vcsAvailable_4;
    R2616 <= T2617;
    R2621 <= T2622;
    validVCs_9_0 <= CMeshDOR_9_io_vcsAvailable_0;
    R2626 <= T2627;
    R2631 <= T2632;
    validVCs_9_1 <= CMeshDOR_9_io_vcsAvailable_1;
    R2636 <= T2637;
    R2641 <= T2642;
    validVCs_9_2 <= CMeshDOR_9_io_vcsAvailable_2;
    R2646 <= T2647;
    R2651 <= T2652;
    validVCs_9_3 <= CMeshDOR_9_io_vcsAvailable_3;
    R2656 <= T2657;
    R2661 <= T2662;
    validVCs_9_4 <= CMeshDOR_9_io_vcsAvailable_4;
    R2666 <= T2667;
    R2671 <= T2672;
    if(reset) begin
      R2675 <= 3'h0;
    end else if(T1670) begin
      R2675 <= T2677;
    end
    if(reset) begin
      R2683 <= 8'h0;
    end else begin
      R2683 <= T2684;
    end
    if(reset) begin
      R2688 <= 1'h1;
    end else begin
      R2688 <= T1692;
    end
    if(reset) begin
      R2689 <= 3'h0;
    end else if(T1526) begin
      R2689 <= T2691;
    end
    if(reset) begin
      R2697 <= 8'h0;
    end else begin
      R2697 <= T2698;
    end
    if(reset) begin
      R2702 <= 1'h1;
    end else begin
      R2702 <= T1548;
    end
    if(reset) begin
      R2703 <= 3'h0;
    end else if(T1382) begin
      R2703 <= T2705;
    end
    if(reset) begin
      R2711 <= 8'h0;
    end else begin
      R2711 <= T2712;
    end
    if(reset) begin
      R2716 <= 1'h1;
    end else begin
      R2716 <= T1404;
    end
    if(reset) begin
      R2717 <= 3'h0;
    end else if(T1238) begin
      R2717 <= T2719;
    end
    if(reset) begin
      R2725 <= 8'h0;
    end else begin
      R2725 <= T2726;
    end
    if(reset) begin
      R2730 <= 1'h1;
    end else begin
      R2730 <= T1260;
    end
    if(reset) begin
      R2731 <= 3'h0;
    end else if(T1094) begin
      R2731 <= T2733;
    end
    if(reset) begin
      R2739 <= 8'h0;
    end else begin
      R2739 <= T2740;
    end
    if(reset) begin
      R2744 <= 1'h1;
    end else begin
      R2744 <= T1116;
    end
    if(reset) begin
      R2745 <= 3'h0;
    end else if(T950) begin
      R2745 <= T2747;
    end
    if(reset) begin
      R2753 <= 8'h0;
    end else begin
      R2753 <= T2754;
    end
    if(reset) begin
      R2758 <= 1'h1;
    end else begin
      R2758 <= T972;
    end
    if(reset) begin
      R2759 <= 3'h0;
    end else if(T806) begin
      R2759 <= T2761;
    end
    if(reset) begin
      R2767 <= 8'h0;
    end else begin
      R2767 <= T2768;
    end
    if(reset) begin
      R2772 <= 1'h1;
    end else begin
      R2772 <= T828;
    end
    if(reset) begin
      R2773 <= 3'h0;
    end else if(T662) begin
      R2773 <= T2775;
    end
    if(reset) begin
      R2781 <= 8'h0;
    end else begin
      R2781 <= T2782;
    end
    if(reset) begin
      R2786 <= 1'h1;
    end else begin
      R2786 <= T684;
    end
    if(reset) begin
      R2787 <= 3'h0;
    end else if(T518) begin
      R2787 <= T2789;
    end
    if(reset) begin
      R2795 <= 8'h0;
    end else begin
      R2795 <= T2796;
    end
    if(reset) begin
      R2800 <= 1'h1;
    end else begin
      R2800 <= T540;
    end
    if(reset) begin
      R2801 <= 3'h0;
    end else if(T374) begin
      R2801 <= T2803;
    end
    if(reset) begin
      R2809 <= 8'h0;
    end else begin
      R2809 <= T2810;
    end
    if(reset) begin
      R2814 <= 1'h1;
    end else begin
      R2814 <= T396;
    end
    R3097 <= T2094;
    if(reset) begin
      R3098 <= T3099;
    end else begin
      R3098 <= switch_io_outPorts_0_x;
    end
    R3100 <= T2031;
    if(reset) begin
      R3101 <= T3102;
    end else begin
      R3101 <= switch_io_outPorts_1_x;
    end
    R3103 <= T1968;
    if(reset) begin
      R3104 <= T3105;
    end else begin
      R3104 <= switch_io_outPorts_2_x;
    end
    R3106 <= T1905;
    if(reset) begin
      R3107 <= T3108;
    end else begin
      R3107 <= switch_io_outPorts_3_x;
    end
    R3109 <= T1722;
    if(reset) begin
      R3110 <= T3111;
    end else begin
      R3110 <= switch_io_outPorts_4_x;
    end
  end
endmodule

module VCRouterWrapper_0(input clk, input reset,
    input [54:0] io_inChannels_4_flit_x,
    input  io_inChannels_4_flitValid,
    output io_inChannels_4_credit_1_grant,
    output io_inChannels_4_credit_0_grant,
    input [54:0] io_inChannels_3_flit_x,
    input  io_inChannels_3_flitValid,
    output io_inChannels_3_credit_1_grant,
    output io_inChannels_3_credit_0_grant,
    input [54:0] io_inChannels_2_flit_x,
    input  io_inChannels_2_flitValid,
    output io_inChannels_2_credit_1_grant,
    output io_inChannels_2_credit_0_grant,
    input [54:0] io_inChannels_1_flit_x,
    input  io_inChannels_1_flitValid,
    output io_inChannels_1_credit_1_grant,
    output io_inChannels_1_credit_0_grant,
    input [54:0] io_inChannels_0_flit_x,
    input  io_inChannels_0_flitValid,
    output io_inChannels_0_credit_1_grant,
    output io_inChannels_0_credit_0_grant,
    output[54:0] io_outChannels_4_flit_x,
    output io_outChannels_4_flitValid,
    input  io_outChannels_4_credit_1_grant,
    input  io_outChannels_4_credit_0_grant,
    output[54:0] io_outChannels_3_flit_x,
    output io_outChannels_3_flitValid,
    input  io_outChannels_3_credit_1_grant,
    input  io_outChannels_3_credit_0_grant,
    output[54:0] io_outChannels_2_flit_x,
    output io_outChannels_2_flitValid,
    input  io_outChannels_2_credit_1_grant,
    input  io_outChannels_2_credit_0_grant,
    output[54:0] io_outChannels_1_flit_x,
    output io_outChannels_1_flitValid,
    input  io_outChannels_1_credit_1_grant,
    input  io_outChannels_1_credit_0_grant,
    output[54:0] io_outChannels_0_flit_x,
    output io_outChannels_0_flitValid,
    input  io_outChannels_0_credit_1_grant,
    input  io_outChannels_0_credit_0_grant,
    output[31:0] io_counters_1_counterVal,
    output[7:0] io_counters_1_counterIndex,
    output[31:0] io_counters_0_counterVal,
    output[7:0] io_counters_0_counterIndex,
    input  io_bypass
);

  wire bp_io_x_inChannels_4_credit_1_grant;
  wire bp_io_x_inChannels_4_credit_0_grant;
  wire bp_io_x_inChannels_3_credit_1_grant;
  wire bp_io_x_inChannels_3_credit_0_grant;
  wire bp_io_x_inChannels_2_credit_1_grant;
  wire bp_io_x_inChannels_2_credit_0_grant;
  wire bp_io_x_inChannels_1_credit_1_grant;
  wire bp_io_x_inChannels_1_credit_0_grant;
  wire bp_io_x_inChannels_0_credit_1_grant;
  wire bp_io_x_inChannels_0_credit_0_grant;
  wire[54:0] bp_io_x_outChannels_4_flit_x;
  wire bp_io_x_outChannels_4_flitValid;
  wire[54:0] bp_io_x_outChannels_3_flit_x;
  wire bp_io_x_outChannels_3_flitValid;
  wire[54:0] bp_io_x_outChannels_2_flit_x;
  wire bp_io_x_outChannels_2_flitValid;
  wire[54:0] bp_io_x_outChannels_1_flit_x;
  wire bp_io_x_outChannels_1_flitValid;
  wire[54:0] bp_io_x_outChannels_0_flit_x;
  wire bp_io_x_outChannels_0_flitValid;
  wire[31:0] bp_io_x_counters_1_counterVal;
  wire[7:0] bp_io_x_counters_1_counterIndex;
  wire[31:0] bp_io_x_counters_0_counterVal;
  wire[7:0] bp_io_x_counters_0_counterIndex;
  wire[54:0] bp_io_y_inChannels_4_flit_x;
  wire bp_io_y_inChannels_4_flitValid;
  wire[54:0] bp_io_y_inChannels_3_flit_x;
  wire bp_io_y_inChannels_3_flitValid;
  wire[54:0] bp_io_y_inChannels_2_flit_x;
  wire bp_io_y_inChannels_2_flitValid;
  wire[54:0] bp_io_y_inChannels_1_flit_x;
  wire bp_io_y_inChannels_1_flitValid;
  wire[54:0] bp_io_y_inChannels_0_flit_x;
  wire bp_io_y_inChannels_0_flitValid;
  wire bp_io_y_outChannels_4_credit_1_grant;
  wire bp_io_y_outChannels_4_credit_0_grant;
  wire bp_io_y_outChannels_3_credit_1_grant;
  wire bp_io_y_outChannels_3_credit_0_grant;
  wire bp_io_y_outChannels_2_credit_1_grant;
  wire bp_io_y_outChannels_2_credit_0_grant;
  wire bp_io_y_outChannels_1_credit_1_grant;
  wire bp_io_y_outChannels_1_credit_0_grant;
  wire bp_io_y_outChannels_0_credit_1_grant;
  wire bp_io_y_outChannels_0_credit_0_grant;
  wire x_io_inChannels_4_credit_1_grant;
  wire x_io_inChannels_4_credit_0_grant;
  wire x_io_inChannels_3_credit_1_grant;
  wire x_io_inChannels_3_credit_0_grant;
  wire x_io_inChannels_2_credit_1_grant;
  wire x_io_inChannels_2_credit_0_grant;
  wire x_io_inChannels_1_credit_1_grant;
  wire x_io_inChannels_1_credit_0_grant;
  wire x_io_inChannels_0_credit_1_grant;
  wire x_io_inChannels_0_credit_0_grant;
  wire[54:0] x_io_outChannels_4_flit_x;
  wire x_io_outChannels_4_flitValid;
  wire[54:0] x_io_outChannels_3_flit_x;
  wire x_io_outChannels_3_flitValid;
  wire[54:0] x_io_outChannels_2_flit_x;
  wire x_io_outChannels_2_flitValid;
  wire[54:0] x_io_outChannels_1_flit_x;
  wire x_io_outChannels_1_flitValid;
  wire[54:0] x_io_outChannels_0_flit_x;
  wire x_io_outChannels_0_flitValid;
  wire[31:0] x_io_counters_0_counterVal;


  assign io_counters_0_counterIndex = bp_io_x_counters_0_counterIndex;
  assign io_counters_0_counterVal = bp_io_x_counters_0_counterVal;
  assign io_counters_1_counterIndex = bp_io_x_counters_1_counterIndex;
  assign io_counters_1_counterVal = bp_io_x_counters_1_counterVal;
  assign io_outChannels_0_flitValid = bp_io_x_outChannels_0_flitValid;
  assign io_outChannels_0_flit_x = bp_io_x_outChannels_0_flit_x;
  assign io_outChannels_1_flitValid = bp_io_x_outChannels_1_flitValid;
  assign io_outChannels_1_flit_x = bp_io_x_outChannels_1_flit_x;
  assign io_outChannels_2_flitValid = bp_io_x_outChannels_2_flitValid;
  assign io_outChannels_2_flit_x = bp_io_x_outChannels_2_flit_x;
  assign io_outChannels_3_flitValid = bp_io_x_outChannels_3_flitValid;
  assign io_outChannels_3_flit_x = bp_io_x_outChannels_3_flit_x;
  assign io_outChannels_4_flitValid = bp_io_x_outChannels_4_flitValid;
  assign io_outChannels_4_flit_x = bp_io_x_outChannels_4_flit_x;
  assign io_inChannels_0_credit_0_grant = bp_io_x_inChannels_0_credit_0_grant;
  assign io_inChannels_0_credit_1_grant = bp_io_x_inChannels_0_credit_1_grant;
  assign io_inChannels_1_credit_0_grant = bp_io_x_inChannels_1_credit_0_grant;
  assign io_inChannels_1_credit_1_grant = bp_io_x_inChannels_1_credit_1_grant;
  assign io_inChannels_2_credit_0_grant = bp_io_x_inChannels_2_credit_0_grant;
  assign io_inChannels_2_credit_1_grant = bp_io_x_inChannels_2_credit_1_grant;
  assign io_inChannels_3_credit_0_grant = bp_io_x_inChannels_3_credit_0_grant;
  assign io_inChannels_3_credit_1_grant = bp_io_x_inChannels_3_credit_1_grant;
  assign io_inChannels_4_credit_0_grant = bp_io_x_inChannels_4_credit_0_grant;
  assign io_inChannels_4_credit_1_grant = bp_io_x_inChannels_4_credit_1_grant;

  wire clkOut;
  VCRouterBypass bp(.clk(clk), .reset(reset),
       .io_x_inChannels_4_flit_x( io_inChannels_4_flit_x ),
       .io_x_inChannels_4_flitValid( io_inChannels_4_flitValid ),
       .io_x_inChannels_4_credit_1_grant( bp_io_x_inChannels_4_credit_1_grant ),
       .io_x_inChannels_4_credit_0_grant( bp_io_x_inChannels_4_credit_0_grant ),
       .io_x_inChannels_3_flit_x( io_inChannels_3_flit_x ),
       .io_x_inChannels_3_flitValid( io_inChannels_3_flitValid ),
       .io_x_inChannels_3_credit_1_grant( bp_io_x_inChannels_3_credit_1_grant ),
       .io_x_inChannels_3_credit_0_grant( bp_io_x_inChannels_3_credit_0_grant ),
       .io_x_inChannels_2_flit_x( io_inChannels_2_flit_x ),
       .io_x_inChannels_2_flitValid( io_inChannels_2_flitValid ),
       .io_x_inChannels_2_credit_1_grant( bp_io_x_inChannels_2_credit_1_grant ),
       .io_x_inChannels_2_credit_0_grant( bp_io_x_inChannels_2_credit_0_grant ),
       .io_x_inChannels_1_flit_x( io_inChannels_1_flit_x ),
       .io_x_inChannels_1_flitValid( io_inChannels_1_flitValid ),
       .io_x_inChannels_1_credit_1_grant( bp_io_x_inChannels_1_credit_1_grant ),
       .io_x_inChannels_1_credit_0_grant( bp_io_x_inChannels_1_credit_0_grant ),
       .io_x_inChannels_0_flit_x( io_inChannels_0_flit_x ),
       .io_x_inChannels_0_flitValid( io_inChannels_0_flitValid ),
       .io_x_inChannels_0_credit_1_grant( bp_io_x_inChannels_0_credit_1_grant ),
       .io_x_inChannels_0_credit_0_grant( bp_io_x_inChannels_0_credit_0_grant ),
       .io_x_outChannels_4_flit_x( bp_io_x_outChannels_4_flit_x ),
       .io_x_outChannels_4_flitValid( bp_io_x_outChannels_4_flitValid ),
       .io_x_outChannels_4_credit_1_grant( io_outChannels_4_credit_1_grant ),
       .io_x_outChannels_4_credit_0_grant( io_outChannels_4_credit_0_grant ),
       .io_x_outChannels_3_flit_x( bp_io_x_outChannels_3_flit_x ),
       .io_x_outChannels_3_flitValid( bp_io_x_outChannels_3_flitValid ),
       .io_x_outChannels_3_credit_1_grant( io_outChannels_3_credit_1_grant ),
       .io_x_outChannels_3_credit_0_grant( io_outChannels_3_credit_0_grant ),
       .io_x_outChannels_2_flit_x( bp_io_x_outChannels_2_flit_x ),
       .io_x_outChannels_2_flitValid( bp_io_x_outChannels_2_flitValid ),
       .io_x_outChannels_2_credit_1_grant( io_outChannels_2_credit_1_grant ),
       .io_x_outChannels_2_credit_0_grant( io_outChannels_2_credit_0_grant ),
       .io_x_outChannels_1_flit_x( bp_io_x_outChannels_1_flit_x ),
       .io_x_outChannels_1_flitValid( bp_io_x_outChannels_1_flitValid ),
       .io_x_outChannels_1_credit_1_grant( io_outChannels_1_credit_1_grant ),
       .io_x_outChannels_1_credit_0_grant( io_outChannels_1_credit_0_grant ),
       .io_x_outChannels_0_flit_x( bp_io_x_outChannels_0_flit_x ),
       .io_x_outChannels_0_flitValid( bp_io_x_outChannels_0_flitValid ),
       .io_x_outChannels_0_credit_1_grant( io_outChannels_0_credit_1_grant ),
       .io_x_outChannels_0_credit_0_grant( io_outChannels_0_credit_0_grant ),
       .io_x_counters_1_counterVal( bp_io_x_counters_1_counterVal ),
       .io_x_counters_1_counterIndex( bp_io_x_counters_1_counterIndex ),
       .io_x_counters_0_counterVal( bp_io_x_counters_0_counterVal ),
       .io_x_counters_0_counterIndex( bp_io_x_counters_0_counterIndex ),
       .io_y_inChannels_4_flit_x( bp_io_y_inChannels_4_flit_x ),
       .io_y_inChannels_4_flitValid( bp_io_y_inChannels_4_flitValid ),
       .io_y_inChannels_4_credit_1_grant( x_io_inChannels_4_credit_1_grant ),
       .io_y_inChannels_4_credit_0_grant( x_io_inChannels_4_credit_0_grant ),
       .io_y_inChannels_3_flit_x( bp_io_y_inChannels_3_flit_x ),
       .io_y_inChannels_3_flitValid( bp_io_y_inChannels_3_flitValid ),
       .io_y_inChannels_3_credit_1_grant( x_io_inChannels_3_credit_1_grant ),
       .io_y_inChannels_3_credit_0_grant( x_io_inChannels_3_credit_0_grant ),
       .io_y_inChannels_2_flit_x( bp_io_y_inChannels_2_flit_x ),
       .io_y_inChannels_2_flitValid( bp_io_y_inChannels_2_flitValid ),
       .io_y_inChannels_2_credit_1_grant( x_io_inChannels_2_credit_1_grant ),
       .io_y_inChannels_2_credit_0_grant( x_io_inChannels_2_credit_0_grant ),
       .io_y_inChannels_1_flit_x( bp_io_y_inChannels_1_flit_x ),
       .io_y_inChannels_1_flitValid( bp_io_y_inChannels_1_flitValid ),
       .io_y_inChannels_1_credit_1_grant( x_io_inChannels_1_credit_1_grant ),
       .io_y_inChannels_1_credit_0_grant( x_io_inChannels_1_credit_0_grant ),
       .io_y_inChannels_0_flit_x( bp_io_y_inChannels_0_flit_x ),
       .io_y_inChannels_0_flitValid( bp_io_y_inChannels_0_flitValid ),
       .io_y_inChannels_0_credit_1_grant( x_io_inChannels_0_credit_1_grant ),
       .io_y_inChannels_0_credit_0_grant( x_io_inChannels_0_credit_0_grant ),
       .io_y_outChannels_4_flit_x( x_io_outChannels_4_flit_x ),
       .io_y_outChannels_4_flitValid( x_io_outChannels_4_flitValid ),
       .io_y_outChannels_4_credit_1_grant( bp_io_y_outChannels_4_credit_1_grant ),
       .io_y_outChannels_4_credit_0_grant( bp_io_y_outChannels_4_credit_0_grant ),
       .io_y_outChannels_3_flit_x( x_io_outChannels_3_flit_x ),
       .io_y_outChannels_3_flitValid( x_io_outChannels_3_flitValid ),
       .io_y_outChannels_3_credit_1_grant( bp_io_y_outChannels_3_credit_1_grant ),
       .io_y_outChannels_3_credit_0_grant( bp_io_y_outChannels_3_credit_0_grant ),
       .io_y_outChannels_2_flit_x( x_io_outChannels_2_flit_x ),
       .io_y_outChannels_2_flitValid( x_io_outChannels_2_flitValid ),
       .io_y_outChannels_2_credit_1_grant( bp_io_y_outChannels_2_credit_1_grant ),
       .io_y_outChannels_2_credit_0_grant( bp_io_y_outChannels_2_credit_0_grant ),
       .io_y_outChannels_1_flit_x( x_io_outChannels_1_flit_x ),
       .io_y_outChannels_1_flitValid( x_io_outChannels_1_flitValid ),
       .io_y_outChannels_1_credit_1_grant( bp_io_y_outChannels_1_credit_1_grant ),
       .io_y_outChannels_1_credit_0_grant( bp_io_y_outChannels_1_credit_0_grant ),
       .io_y_outChannels_0_flit_x( x_io_outChannels_0_flit_x ),
       .io_y_outChannels_0_flitValid( x_io_outChannels_0_flitValid ),
       .io_y_outChannels_0_credit_1_grant( bp_io_y_outChannels_0_credit_1_grant ),
       .io_y_outChannels_0_credit_0_grant( bp_io_y_outChannels_0_credit_0_grant ),
       //.io_y_counters_1_counterVal(  )
       //.io_y_counters_1_counterIndex(  )
       .io_y_counters_0_counterVal( x_io_counters_0_counterVal ),
       //.io_y_counters_0_counterIndex(  )
       .io_bypass( io_bypass ),
       .io_clkOut(clkOut)
  );
  SimpleVCRouter_0 x(.clk(clkOut), .reset(reset),
       .io_inChannels_4_flit_x( bp_io_y_inChannels_4_flit_x ),
       .io_inChannels_4_flitValid( bp_io_y_inChannels_4_flitValid ),
       .io_inChannels_4_credit_1_grant( x_io_inChannels_4_credit_1_grant ),
       .io_inChannels_4_credit_0_grant( x_io_inChannels_4_credit_0_grant ),
       .io_inChannels_3_flit_x( bp_io_y_inChannels_3_flit_x ),
       .io_inChannels_3_flitValid( bp_io_y_inChannels_3_flitValid ),
       .io_inChannels_3_credit_1_grant( x_io_inChannels_3_credit_1_grant ),
       .io_inChannels_3_credit_0_grant( x_io_inChannels_3_credit_0_grant ),
       .io_inChannels_2_flit_x( bp_io_y_inChannels_2_flit_x ),
       .io_inChannels_2_flitValid( bp_io_y_inChannels_2_flitValid ),
       .io_inChannels_2_credit_1_grant( x_io_inChannels_2_credit_1_grant ),
       .io_inChannels_2_credit_0_grant( x_io_inChannels_2_credit_0_grant ),
       .io_inChannels_1_flit_x( bp_io_y_inChannels_1_flit_x ),
       .io_inChannels_1_flitValid( bp_io_y_inChannels_1_flitValid ),
       .io_inChannels_1_credit_1_grant( x_io_inChannels_1_credit_1_grant ),
       .io_inChannels_1_credit_0_grant( x_io_inChannels_1_credit_0_grant ),
       .io_inChannels_0_flit_x( bp_io_y_inChannels_0_flit_x ),
       .io_inChannels_0_flitValid( bp_io_y_inChannels_0_flitValid ),
       .io_inChannels_0_credit_1_grant( x_io_inChannels_0_credit_1_grant ),
       .io_inChannels_0_credit_0_grant( x_io_inChannels_0_credit_0_grant ),
       .io_outChannels_4_flit_x( x_io_outChannels_4_flit_x ),
       .io_outChannels_4_flitValid( x_io_outChannels_4_flitValid ),
       .io_outChannels_4_credit_1_grant( bp_io_y_outChannels_4_credit_1_grant ),
       .io_outChannels_4_credit_0_grant( bp_io_y_outChannels_4_credit_0_grant ),
       .io_outChannels_3_flit_x( x_io_outChannels_3_flit_x ),
       .io_outChannels_3_flitValid( x_io_outChannels_3_flitValid ),
       .io_outChannels_3_credit_1_grant( bp_io_y_outChannels_3_credit_1_grant ),
       .io_outChannels_3_credit_0_grant( bp_io_y_outChannels_3_credit_0_grant ),
       .io_outChannels_2_flit_x( x_io_outChannels_2_flit_x ),
       .io_outChannels_2_flitValid( x_io_outChannels_2_flitValid ),
       .io_outChannels_2_credit_1_grant( bp_io_y_outChannels_2_credit_1_grant ),
       .io_outChannels_2_credit_0_grant( bp_io_y_outChannels_2_credit_0_grant ),
       .io_outChannels_1_flit_x( x_io_outChannels_1_flit_x ),
       .io_outChannels_1_flitValid( x_io_outChannels_1_flitValid ),
       .io_outChannels_1_credit_1_grant( bp_io_y_outChannels_1_credit_1_grant ),
       .io_outChannels_1_credit_0_grant( bp_io_y_outChannels_1_credit_0_grant ),
       .io_outChannels_0_flit_x( x_io_outChannels_0_flit_x ),
       .io_outChannels_0_flitValid( x_io_outChannels_0_flitValid ),
       .io_outChannels_0_credit_1_grant( bp_io_y_outChannels_0_credit_1_grant ),
       .io_outChannels_0_credit_0_grant( bp_io_y_outChannels_0_credit_0_grant ),
       //.io_counters_1_counterVal(  )
       //.io_counters_1_counterIndex(  )
       .io_counters_0_counterVal( x_io_counters_0_counterVal )
       //.io_counters_0_counterIndex(  )
       //.io_bypass(  )
  );
endmodule

module BusProbe_0(input clk, input reset,
    //input [54:0] io_inFlit_4_x
    //input [54:0] io_inFlit_3_x
    //input [54:0] io_inFlit_2_x
    input [54:0] io_inFlit_1_x,
    //input [54:0] io_inFlit_0_x
    input  io_inValid_4,
    input  io_inValid_3,
    input  io_inValid_2,
    input  io_inValid_1,
    input  io_inValid_0,
    input  io_routerCord,
    //input  io_startRecording
    output[15:0] io_cyclesChannelBusy_4,
    output[15:0] io_cyclesChannelBusy_3,
    output[15:0] io_cyclesChannelBusy_2,
    output[15:0] io_cyclesChannelBusy_1,
    output[15:0] io_cyclesChannelBusy_0,
    output[15:0] io_cyclesRouterBusy
);

  reg[0:0] T0;
  reg [15:0] cyclesRouterBusy;
  wire[15:0] T29;
  wire[15:0] T1;
  wire[15:0] T2;
  wire T3;
  wire[4:0] T4;
  wire[4:0] T5;
  wire[2:0] T6;
  wire[1:0] T7;
  reg  cyclesChannelBusyScoreboard_0;
  wire T30;
  wire T8;
  wire T9;
  reg  cyclesChannelBusyScoreboard_1;
  wire T31;
  wire T10;
  wire T11;
  reg  cyclesChannelBusyScoreboard_2;
  wire T32;
  wire T12;
  wire T13;
  wire[1:0] T14;
  reg  cyclesChannelBusyScoreboard_3;
  wire T33;
  wire T15;
  wire T16;
  reg  cyclesChannelBusyScoreboard_4;
  wire T34;
  wire T17;
  wire T18;
  reg [15:0] cyclesChannelBusy_0;
  wire[15:0] T35;
  wire[15:0] T19;
  wire[15:0] T20;
  reg [15:0] cyclesChannelBusy_1;
  wire[15:0] T36;
  wire[15:0] T21;
  wire[15:0] T22;
  reg [15:0] cyclesChannelBusy_2;
  wire[15:0] T37;
  wire[15:0] T23;
  wire[15:0] T24;
  reg [15:0] cyclesChannelBusy_3;
  wire[15:0] T38;
  wire[15:0] T25;
  wire[15:0] T26;
  reg [15:0] cyclesChannelBusy_4;
  wire[15:0] T39;
  wire[15:0] T27;
  wire[15:0] T28;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    T0 = 1'b0;
    cyclesRouterBusy = {1{1'b0}};
    cyclesChannelBusyScoreboard_0 = {1{1'b0}};
    cyclesChannelBusyScoreboard_1 = {1{1'b0}};
    cyclesChannelBusyScoreboard_2 = {1{1'b0}};
    cyclesChannelBusyScoreboard_3 = {1{1'b0}};
    cyclesChannelBusyScoreboard_4 = {1{1'b0}};
    cyclesChannelBusy_0 = {1{1'b0}};
    cyclesChannelBusy_1 = {1{1'b0}};
    cyclesChannelBusy_2 = {1{1'b0}};
    cyclesChannelBusy_3 = {1{1'b0}};
    cyclesChannelBusy_4 = {1{1'b0}};
  end
// synthesis translate_on
`endif

  assign io_cyclesRouterBusy = cyclesRouterBusy;
  assign T29 = reset ? 16'h0 : T1;
  assign T1 = T3 ? T2 : cyclesRouterBusy;
  assign T2 = cyclesRouterBusy + 16'h1;
  assign T3 = T4 != 5'h0;
  assign T4 = T5;
  assign T5 = {T14, T6};
  assign T6 = {cyclesChannelBusyScoreboard_2, T7};
  assign T7 = {cyclesChannelBusyScoreboard_1, cyclesChannelBusyScoreboard_0};
  assign T30 = reset ? 1'h0 : T8;
  assign T8 = T9 == 1'h0;
  assign T9 = io_inValid_0 ^ 1'h1;
  assign T31 = reset ? 1'h0 : T10;
  assign T10 = T11 == 1'h0;
  assign T11 = io_inValid_1 ^ 1'h1;
  assign T32 = reset ? 1'h0 : T12;
  assign T12 = T13 == 1'h0;
  assign T13 = io_inValid_2 ^ 1'h1;
  assign T14 = {cyclesChannelBusyScoreboard_4, cyclesChannelBusyScoreboard_3};
  assign T33 = reset ? 1'h0 : T15;
  assign T15 = T16 == 1'h0;
  assign T16 = io_inValid_3 ^ 1'h1;
  assign T34 = reset ? 1'h0 : T17;
  assign T17 = T18 == 1'h0;
  assign T18 = io_inValid_4 ^ 1'h1;
  assign io_cyclesChannelBusy_0 = cyclesChannelBusy_0;
  assign T35 = reset ? 16'h0 : T19;
  assign T19 = io_inValid_0 ? T20 : cyclesChannelBusy_0;
  assign T20 = cyclesChannelBusy_0 + 16'h1;
  assign io_cyclesChannelBusy_1 = cyclesChannelBusy_1;
  assign T36 = reset ? 16'h0 : T21;
  assign T21 = io_inValid_1 ? T22 : cyclesChannelBusy_1;
  assign T22 = cyclesChannelBusy_1 + 16'h1;
  assign io_cyclesChannelBusy_2 = cyclesChannelBusy_2;
  assign T37 = reset ? 16'h0 : T23;
  assign T23 = io_inValid_2 ? T24 : cyclesChannelBusy_2;
  assign T24 = cyclesChannelBusy_2 + 16'h1;
  assign io_cyclesChannelBusy_3 = cyclesChannelBusy_3;
  assign T38 = reset ? 16'h0 : T25;
  assign T25 = io_inValid_3 ? T26 : cyclesChannelBusy_3;
  assign T26 = cyclesChannelBusy_3 + 16'h1;
  assign io_cyclesChannelBusy_4 = cyclesChannelBusy_4;
  assign T39 = reset ? 16'h0 : T27;
  assign T27 = io_inValid_4 ? T28 : cyclesChannelBusy_4;
  assign T28 = cyclesChannelBusy_4 + 16'h1;

  always @(posedge clk) begin
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T0 <= 1'b1;
  if(!1'h1 && T0 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "BusProbe: RouterRadix must be > 1");
    $finish;
  end
// synthesis translate_on
`endif
    if(reset) begin
      cyclesRouterBusy <= 16'h0;
    end else if(T3) begin
      cyclesRouterBusy <= T2;
    end
    if(reset) begin
      cyclesChannelBusyScoreboard_0 <= 1'h0;
    end else begin
      cyclesChannelBusyScoreboard_0 <= T8;
    end
    if(reset) begin
      cyclesChannelBusyScoreboard_1 <= 1'h0;
    end else begin
      cyclesChannelBusyScoreboard_1 <= T10;
    end
    if(reset) begin
      cyclesChannelBusyScoreboard_2 <= 1'h0;
    end else begin
      cyclesChannelBusyScoreboard_2 <= T12;
    end
    if(reset) begin
      cyclesChannelBusyScoreboard_3 <= 1'h0;
    end else begin
      cyclesChannelBusyScoreboard_3 <= T15;
    end
    if(reset) begin
      cyclesChannelBusyScoreboard_4 <= 1'h0;
    end else begin
      cyclesChannelBusyScoreboard_4 <= T17;
    end
    if(reset) begin
      cyclesChannelBusy_0 <= 16'h0;
    end else if(io_inValid_0) begin
      cyclesChannelBusy_0 <= T20;
    end
    if(reset) begin
      cyclesChannelBusy_1 <= 16'h0;
    end else if(io_inValid_1) begin
      cyclesChannelBusy_1 <= T22;
    end
    if(reset) begin
      cyclesChannelBusy_2 <= 16'h0;
    end else if(io_inValid_2) begin
      cyclesChannelBusy_2 <= T24;
    end
    if(reset) begin
      cyclesChannelBusy_3 <= 16'h0;
    end else if(io_inValid_3) begin
      cyclesChannelBusy_3 <= T26;
    end
    if(reset) begin
      cyclesChannelBusy_4 <= 16'h0;
    end else if(io_inValid_4) begin
      cyclesChannelBusy_4 <= T28;
    end
  end
endmodule

module CreditBuffer(input clk, input reset,
    input [54:0] io_in_4_flit_x,
    input  io_in_4_flitValid,
    output io_in_4_credit_1_grant,
    output io_in_4_credit_0_grant,
    input [54:0] io_in_3_flit_x,
    input  io_in_3_flitValid,
    output io_in_3_credit_1_grant,
    output io_in_3_credit_0_grant,
    input [54:0] io_in_2_flit_x,
    input  io_in_2_flitValid,
    output io_in_2_credit_1_grant,
    output io_in_2_credit_0_grant,
    input [54:0] io_in_1_flit_x,
    input  io_in_1_flitValid,
    output io_in_1_credit_1_grant,
    output io_in_1_credit_0_grant,
    input [54:0] io_in_0_flit_x,
    input  io_in_0_flitValid,
    output io_in_0_credit_1_grant,
    output io_in_0_credit_0_grant,
    output[54:0] io_out_4_flit_x,
    output io_out_4_flitValid,
    input  io_out_4_credit_1_grant,
    input  io_out_4_credit_0_grant,
    output[54:0] io_out_3_flit_x,
    output io_out_3_flitValid,
    input  io_out_3_credit_1_grant,
    input  io_out_3_credit_0_grant,
    output[54:0] io_out_2_flit_x,
    output io_out_2_flitValid,
    input  io_out_2_credit_1_grant,
    input  io_out_2_credit_0_grant,
    output[54:0] io_out_1_flit_x,
    output io_out_1_flitValid,
    input  io_out_1_credit_1_grant,
    input  io_out_1_credit_0_grant,
    output[54:0] io_out_0_flit_x,
    output io_out_0_flitValid,
    input  io_out_0_credit_1_grant,
    input  io_out_0_credit_0_grant
);

  wire T0;
  reg  R1;
  wire T20;
  wire T2;
  reg  R3;
  wire T21;
  wire T4;
  reg  R5;
  wire T22;
  wire T6;
  reg  R7;
  wire T23;
  wire T8;
  reg  R9;
  wire T24;
  wire T10;
  reg  R11;
  wire T25;
  wire T12;
  reg  R13;
  wire T26;
  wire T14;
  reg  R15;
  wire T27;
  wire T16;
  reg  R17;
  wire T28;
  wire T18;
  reg  R19;
  wire T29;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    R1 = {1{1'b0}};
    R3 = {1{1'b0}};
    R5 = {1{1'b0}};
    R7 = {1{1'b0}};
    R9 = {1{1'b0}};
    R11 = {1{1'b0}};
    R13 = {1{1'b0}};
    R15 = {1{1'b0}};
    R17 = {1{1'b0}};
    R19 = {1{1'b0}};
  end
// synthesis translate_on
`endif

  assign io_out_0_flitValid = io_in_0_flitValid;
  assign io_out_0_flit_x = io_in_0_flit_x;
  assign io_out_1_flitValid = io_in_1_flitValid;
  assign io_out_1_flit_x = io_in_1_flit_x;
  assign io_out_2_flitValid = io_in_2_flitValid;
  assign io_out_2_flit_x = io_in_2_flit_x;
  assign io_out_3_flitValid = io_in_3_flitValid;
  assign io_out_3_flit_x = io_in_3_flit_x;
  assign io_out_4_flitValid = io_in_4_flitValid;
  assign io_out_4_flit_x = io_in_4_flit_x;
  assign io_in_0_credit_0_grant = T0;
  assign T0 = R1;
  assign T20 = reset ? 1'h0 : io_out_0_credit_0_grant;
  assign io_in_0_credit_1_grant = T2;
  assign T2 = R3;
  assign T21 = reset ? 1'h0 : io_out_0_credit_1_grant;
  assign io_in_1_credit_0_grant = T4;
  assign T4 = R5;
  assign T22 = reset ? 1'h0 : io_out_1_credit_0_grant;
  assign io_in_1_credit_1_grant = T6;
  assign T6 = R7;
  assign T23 = reset ? 1'h0 : io_out_1_credit_1_grant;
  assign io_in_2_credit_0_grant = T8;
  assign T8 = R9;
  assign T24 = reset ? 1'h0 : io_out_2_credit_0_grant;
  assign io_in_2_credit_1_grant = T10;
  assign T10 = R11;
  assign T25 = reset ? 1'h0 : io_out_2_credit_1_grant;
  assign io_in_3_credit_0_grant = T12;
  assign T12 = R13;
  assign T26 = reset ? 1'h0 : io_out_3_credit_0_grant;
  assign io_in_3_credit_1_grant = T14;
  assign T14 = R15;
  assign T27 = reset ? 1'h0 : io_out_3_credit_1_grant;
  assign io_in_4_credit_0_grant = T16;
  assign T16 = R17;
  assign T28 = reset ? 1'h0 : io_out_4_credit_0_grant;
  assign io_in_4_credit_1_grant = T18;
  assign T18 = R19;
  assign T29 = reset ? 1'h0 : io_out_4_credit_1_grant;

  always @(posedge clk) begin
    if(reset) begin
      R1 <= 1'h0;
    end else begin
      R1 <= io_out_0_credit_0_grant;
    end
    if(reset) begin
      R3 <= 1'h0;
    end else begin
      R3 <= io_out_0_credit_1_grant;
    end
    if(reset) begin
      R5 <= 1'h0;
    end else begin
      R5 <= io_out_1_credit_0_grant;
    end
    if(reset) begin
      R7 <= 1'h0;
    end else begin
      R7 <= io_out_1_credit_1_grant;
    end
    if(reset) begin
      R9 <= 1'h0;
    end else begin
      R9 <= io_out_2_credit_0_grant;
    end
    if(reset) begin
      R11 <= 1'h0;
    end else begin
      R11 <= io_out_2_credit_1_grant;
    end
    if(reset) begin
      R13 <= 1'h0;
    end else begin
      R13 <= io_out_3_credit_0_grant;
    end
    if(reset) begin
      R15 <= 1'h0;
    end else begin
      R15 <= io_out_3_credit_1_grant;
    end
    if(reset) begin
      R17 <= 1'h0;
    end else begin
      R17 <= io_out_4_credit_0_grant;
    end
    if(reset) begin
      R19 <= 1'h0;
    end else begin
      R19 <= io_out_4_credit_1_grant;
    end
  end
endmodule

module CMeshDOR_1(
    input [15:0] io_inHeadFlit_packetID,
    input  io_inHeadFlit_isTail,
    input  io_inHeadFlit_vcPort,
    input [3:0] io_inHeadFlit_packetType,
    input [1:0] io_inHeadFlit_destination_2,
    input [1:0] io_inHeadFlit_destination_1,
    input [1:0] io_inHeadFlit_destination_0,
    input [2:0] io_inHeadFlit_priorityLevel,
    output[15:0] io_outHeadFlit_packetID,
    output io_outHeadFlit_isTail,
    output io_outHeadFlit_vcPort,
    output[3:0] io_outHeadFlit_packetType,
    output[1:0] io_outHeadFlit_destination_2,
    output[1:0] io_outHeadFlit_destination_1,
    output[1:0] io_outHeadFlit_destination_0,
    output[2:0] io_outHeadFlit_priorityLevel,
    output[2:0] io_result,
    output[1:0] io_vcsAvailable_4,
    output[1:0] io_vcsAvailable_3,
    output[1:0] io_vcsAvailable_2,
    output[1:0] io_vcsAvailable_1,
    output[1:0] io_vcsAvailable_0
);

  wire[1:0] T0;
  wire[1:0] T26;
  wire T1;
  wire[1:0] T2;
  wire[1:0] T27;
  wire T3;
  wire[1:0] T4;
  wire[1:0] T28;
  wire T5;
  wire[1:0] T6;
  wire[1:0] T29;
  wire T7;
  wire[1:0] T8;
  wire[1:0] T30;
  wire T9;
  wire[2:0] T10;
  wire[2:0] resultReduction;
  wire[2:0] T11;
  wire[2:0] dimResults_1;
  wire[2:0] T12;
  wire[2:0] T31;
  wire[1:0] T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire[2:0] dimResults_0;
  wire[2:0] T32;
  wire[1:0] T18;
  wire[1:0] T33;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire[2:0] T34;
  wire T25;


  assign io_vcsAvailable_0 = T0;
  assign T0 = 2'h0 - T26;
  assign T26 = {1'h0, T1};
  assign T1 = io_result == 3'h0;
  assign io_vcsAvailable_1 = T2;
  assign T2 = 2'h0 - T27;
  assign T27 = {1'h0, T3};
  assign T3 = io_result == 3'h1;
  assign io_vcsAvailable_2 = T4;
  assign T4 = 2'h0 - T28;
  assign T28 = {1'h0, T5};
  assign T5 = io_result == 3'h2;
  assign io_vcsAvailable_3 = T6;
  assign T6 = 2'h0 - T29;
  assign T29 = {1'h0, T7};
  assign T7 = io_result == 3'h3;
  assign io_vcsAvailable_4 = T8;
  assign T8 = 2'h0 - T30;
  assign T30 = {1'h0, T9};
  assign T9 = io_result == 3'h4;
  assign io_result = T10;
  assign T10 = T25 ? T34 : resultReduction;
  assign resultReduction = T11;
  assign T11 = T24 ? dimResults_0 : dimResults_1;
  assign dimResults_1 = T12;
  assign T12 = T15 ? 3'h4 : T31;
  assign T31 = {1'h0, T13};
  assign T13 = T14 ? 2'h3 : 2'h0;
  assign T14 = 2'h0 < io_inHeadFlit_destination_1;
  assign T15 = T17 & T16;
  assign T16 = io_inHeadFlit_destination_1 < 2'h0;
  assign T17 = T14 ^ 1'h1;
  assign dimResults_0 = T32;
  assign T32 = {1'h0, T18};
  assign T18 = T21 ? 2'h2 : T33;
  assign T33 = {1'h0, T19};
  assign T19 = T20 ? 1'h1 : 1'h0;
  assign T20 = 2'h1 < io_inHeadFlit_destination_0;
  assign T21 = T23 & T22;
  assign T22 = io_inHeadFlit_destination_0 < 2'h1;
  assign T23 = T20 ^ 1'h1;
  assign T24 = dimResults_0 != 3'h0;
  assign T34 = {1'h0, io_inHeadFlit_destination_2};
  assign T25 = resultReduction == 3'h0;
  assign io_outHeadFlit_priorityLevel = io_inHeadFlit_priorityLevel;
  assign io_outHeadFlit_destination_0 = io_inHeadFlit_destination_0;
  assign io_outHeadFlit_destination_1 = io_inHeadFlit_destination_1;
  assign io_outHeadFlit_destination_2 = io_inHeadFlit_destination_2;
  assign io_outHeadFlit_packetType = io_inHeadFlit_packetType;
  assign io_outHeadFlit_vcPort = io_inHeadFlit_vcPort;
  assign io_outHeadFlit_isTail = io_inHeadFlit_isTail;
  assign io_outHeadFlit_packetID = io_inHeadFlit_packetID;
endmodule

module SimpleVCRouter_1((* gated_clock = "true" *) input clk, input reset,
    input [54:0] io_inChannels_4_flit_x,
    input  io_inChannels_4_flitValid,
    output io_inChannels_4_credit_1_grant,
    output io_inChannels_4_credit_0_grant,
    input [54:0] io_inChannels_3_flit_x,
    input  io_inChannels_3_flitValid,
    output io_inChannels_3_credit_1_grant,
    output io_inChannels_3_credit_0_grant,
    input [54:0] io_inChannels_2_flit_x,
    input  io_inChannels_2_flitValid,
    output io_inChannels_2_credit_1_grant,
    output io_inChannels_2_credit_0_grant,
    input [54:0] io_inChannels_1_flit_x,
    input  io_inChannels_1_flitValid,
    output io_inChannels_1_credit_1_grant,
    output io_inChannels_1_credit_0_grant,
    input [54:0] io_inChannels_0_flit_x,
    input  io_inChannels_0_flitValid,
    output io_inChannels_0_credit_1_grant,
    output io_inChannels_0_credit_0_grant,
    output[54:0] io_outChannels_4_flit_x,
    output io_outChannels_4_flitValid,
    input  io_outChannels_4_credit_1_grant,
    input  io_outChannels_4_credit_0_grant,
    output[54:0] io_outChannels_3_flit_x,
    output io_outChannels_3_flitValid,
    input  io_outChannels_3_credit_1_grant,
    input  io_outChannels_3_credit_0_grant,
    output[54:0] io_outChannels_2_flit_x,
    output io_outChannels_2_flitValid,
    input  io_outChannels_2_credit_1_grant,
    input  io_outChannels_2_credit_0_grant,
    output[54:0] io_outChannels_1_flit_x,
    output io_outChannels_1_flitValid,
    input  io_outChannels_1_credit_1_grant,
    input  io_outChannels_1_credit_0_grant,
    output[54:0] io_outChannels_0_flit_x,
    output io_outChannels_0_flitValid,
    input  io_outChannels_0_credit_1_grant,
    input  io_outChannels_0_credit_0_grant,
    //output[31:0] io_counters_1_counterVal
    //output[7:0] io_counters_1_counterIndex
    output[31:0] io_counters_0_counterVal
    //output[7:0] io_counters_0_counterIndex
    //input  io_bypass
);

  reg[0:0] T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  wire[53:0] T8;
  wire T9;
  wire[30:0] T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  reg[0:0] T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  reg[0:0] T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire[53:0] T30;
  wire T31;
  wire[30:0] T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  reg[0:0] T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  reg[0:0] T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire[53:0] T52;
  wire T53;
  wire[30:0] T54;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  reg[0:0] T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  reg[0:0] T66;
  wire T67;
  wire T68;
  wire T69;
  wire T70;
  wire T71;
  wire T72;
  wire T73;
  wire[53:0] T74;
  wire T75;
  wire[30:0] T76;
  wire T77;
  wire T78;
  wire T79;
  wire T80;
  wire T81;
  wire T82;
  reg[0:0] T83;
  wire T84;
  wire T85;
  wire T86;
  wire T87;
  reg[0:0] T88;
  wire T89;
  wire T90;
  wire T91;
  wire T92;
  wire T93;
  wire T94;
  wire T95;
  wire[53:0] T96;
  wire T97;
  wire[30:0] T98;
  wire T99;
  wire T100;
  wire T101;
  wire T102;
  wire T103;
  wire T104;
  reg[0:0] T105;
  wire T106;
  wire T107;
  wire T108;
  wire T109;
  reg[0:0] T110;
  wire T111;
  wire T112;
  wire T113;
  wire T114;
  wire T115;
  wire T116;
  wire T117;
  wire[53:0] T118;
  wire T119;
  wire[30:0] T120;
  wire T121;
  wire T122;
  wire T123;
  wire T124;
  wire T125;
  wire T126;
  reg[0:0] T127;
  wire T128;
  wire T129;
  wire T130;
  wire T131;
  reg[0:0] T132;
  wire T133;
  wire T134;
  wire T135;
  wire T136;
  wire T137;
  wire T138;
  wire T139;
  wire[53:0] T140;
  wire T141;
  wire[30:0] T142;
  wire T143;
  wire T144;
  wire T145;
  wire T146;
  wire T147;
  wire T148;
  reg[0:0] T149;
  wire T150;
  wire T151;
  wire T152;
  wire T153;
  reg[0:0] T154;
  wire T155;
  wire T156;
  wire T157;
  wire T158;
  wire T159;
  wire T160;
  wire T161;
  wire[53:0] T162;
  wire T163;
  wire[30:0] T164;
  wire T165;
  wire T166;
  wire T167;
  wire T168;
  wire T169;
  wire T170;
  reg[0:0] T171;
  wire T172;
  wire T173;
  wire T174;
  wire T175;
  reg[0:0] T176;
  wire T177;
  wire T178;
  wire T179;
  wire T180;
  wire T181;
  wire T182;
  wire T183;
  wire[53:0] T184;
  wire T185;
  wire[30:0] T186;
  wire T187;
  wire T188;
  wire T189;
  wire T190;
  wire T191;
  wire T192;
  reg[0:0] T193;
  wire T194;
  wire T195;
  wire T196;
  wire T197;
  reg[0:0] T198;
  wire T199;
  wire T200;
  wire T201;
  wire T202;
  wire T203;
  wire T204;
  wire T205;
  wire[53:0] T206;
  wire T207;
  wire[30:0] T208;
  wire T209;
  wire T210;
  wire T211;
  wire T212;
  wire T213;
  wire T214;
  reg[0:0] T215;
  wire T216;
  wire T217;
  wire T218;
  wire T219;
  wire T220;
  wire T221;
  wire T222;
  wire T223;
  wire T224;
  wire[53:0] T225;
  wire T226;
  wire[30:0] T227;
  wire T228;
  wire T229;
  wire T230;
  wire T231;
  wire T232;
  wire T233;
  wire T234;
  wire T235;
  wire T236;
  wire[53:0] T237;
  wire T238;
  wire[30:0] T239;
  wire T240;
  wire T241;
  wire T242;
  wire T243;
  wire T244;
  wire T245;
  wire T246;
  wire T247;
  wire T248;
  wire[53:0] T249;
  wire T250;
  wire[30:0] T251;
  wire T252;
  wire T253;
  wire T254;
  wire T255;
  wire T256;
  wire T257;
  wire T258;
  wire T259;
  wire T260;
  wire[53:0] T261;
  wire T262;
  wire[30:0] T263;
  wire T264;
  wire T265;
  wire T266;
  wire T267;
  wire T268;
  wire T269;
  wire T270;
  wire T271;
  wire T272;
  wire[53:0] T273;
  wire T274;
  wire[30:0] T275;
  wire T276;
  wire T277;
  wire T278;
  wire T279;
  wire[54:0] T280;
  wire[54:0] T281;
  wire T3112;
  reg [54:0] R282;
  wire[54:0] T3113;
  wire[54:0] T283;
  wire[54:0] T3114;
  wire T284;
  wire T285;
  wire[54:0] T286;
  wire[54:0] T287;
  wire T288;
  wire T289;
  wire[1:0] T290;
  wire[1:0] T291;
  wire[1:0] T292;
  wire T293;
  wire[2:0] T294;
  reg [2:0] R295;
  wire[2:0] T3115;
  wire[1:0] T296;
  wire T297;
  wire T298;
  wire T299;
  wire T300;
  wire T301;
  wire T302;
  wire T303;
  wire T304;
  wire creditConsReady_0_0;
  wire creditConsReady_1_0;
  wire T305;
  wire[2:0] T306;
  wire T307;
  wire creditConsReady_2_0;
  wire creditConsReady_3_0;
  wire T308;
  wire T309;
  wire creditConsReady_4_0;
  wire T310;
  wire T311;
  wire T312;
  wire T313;
  wire creditConsReady_0_1;
  wire creditConsReady_1_1;
  wire T314;
  wire T315;
  wire creditConsReady_2_1;
  wire creditConsReady_3_1;
  wire T316;
  wire T317;
  wire creditConsReady_4_1;
  wire T318;
  wire T319;
  wire T3116;
  wire T320;
  wire T321;
  wire[3:0] T322;
  wire[3:0] T323;
  wire[3:0] T324;
  wire T325;
  wire[2:0] T326;
  wire[3:0] T327;
  wire T328;
  wire T329;
  wire T330;
  wire T331;
  wire T332;
  wire T333;
  wire T334;
  wire[2:0] T335;
  wire T336;
  wire T337;
  wire T338;
  wire T339;
  wire T340;
  wire T341;
  wire T342;
  wire T343;
  wire[53:0] T344;
  wire T345;
  wire[30:0] T346;
  wire T347;
  wire T348;
  reg  R349;
  wire T3117;
  wire[2:0] T350;
  wire[30:0] T351;
  wire[54:0] T352;
  wire[1:0] T353;
  wire[1:0] T354;
  wire[1:0] T355;
  wire[3:0] T356;
  wire T357;
  wire T358;
  wire[15:0] T359;
  wire T360;
  wire T361;
  wire T362;
  wire T363;
  wire T364;
  wire T365;
  wire T366;
  wire T367;
  wire T368;
  wire T369;
  wire T370;
  wire T371;
  wire T372;
  wire T373;
  wire T374;
  wire T375;
  wire T376;
  wire T377;
  wire T378;
  wire T379;
  wire T380;
  wire T381;
  wire T382;
  wire T383;
  wire T384;
  wire T385;
  wire T386;
  wire T387;
  wire[54:0] T3118;
  wire[30:0] T388;
  wire[30:0] T389;
  wire[8:0] T390;
  wire[4:0] T391;
  wire[3:0] T392;
  wire[21:0] T393;
  wire[4:0] T394;
  wire[16:0] T395;
  wire T396;
  wire T397;
  wire T398;
  wire T399;
  wire flitsAreTail_9;
  wire T400;
  wire T401;
  wire T402;
  wire T403;
  wire[53:0] T404;
  wire T405;
  wire[30:0] T406;
  wire T407;
  wire T408;
  wire T409;
  wire T410;
  wire T411;
  wire[54:0] T412;
  wire[54:0] T413;
  wire T414;
  wire T415;
  wire T416;
  wire T417;
  wire T418;
  wire T419;
  wire T420;
  wire T421;
  wire T422;
  wire T423;
  wire[54:0] T424;
  wire[54:0] T425;
  wire T3119;
  reg [54:0] R426;
  wire[54:0] T3120;
  wire[54:0] T427;
  wire[54:0] T3121;
  wire T428;
  wire T429;
  wire[54:0] T430;
  wire[54:0] T431;
  wire T432;
  wire T433;
  wire[1:0] T434;
  wire[1:0] T435;
  wire[1:0] T436;
  wire T437;
  wire[2:0] T438;
  reg [2:0] R439;
  wire[2:0] T3122;
  wire[1:0] T440;
  wire T441;
  wire T442;
  wire T443;
  wire T444;
  wire T445;
  wire T446;
  wire T447;
  wire T448;
  wire T449;
  wire[2:0] T450;
  wire T451;
  wire T452;
  wire T453;
  wire T454;
  wire T455;
  wire T456;
  wire T457;
  wire T458;
  wire T459;
  wire T460;
  wire T461;
  wire T462;
  wire T463;
  wire T3123;
  wire T464;
  wire T465;
  wire[3:0] T466;
  wire[3:0] T467;
  wire[3:0] T468;
  wire T469;
  wire[2:0] T470;
  wire[3:0] T471;
  wire T472;
  wire T473;
  wire T474;
  wire T475;
  wire T476;
  wire T477;
  wire T478;
  wire[2:0] T479;
  wire T480;
  wire T481;
  wire T482;
  wire T483;
  wire T484;
  wire T485;
  wire T486;
  wire T487;
  wire[53:0] T488;
  wire T489;
  wire[30:0] T490;
  wire T491;
  wire T492;
  reg  R493;
  wire T3124;
  wire[2:0] T494;
  wire[30:0] T495;
  wire[54:0] T496;
  wire[1:0] T497;
  wire[1:0] T498;
  wire[1:0] T499;
  wire[3:0] T500;
  wire T501;
  wire T502;
  wire[15:0] T503;
  wire T504;
  wire T505;
  wire T506;
  wire T507;
  wire T508;
  wire T509;
  wire T510;
  wire T511;
  wire T512;
  wire T513;
  wire T514;
  wire T515;
  wire T516;
  wire T517;
  wire T518;
  wire T519;
  wire T520;
  wire T521;
  wire T522;
  wire T523;
  wire T524;
  wire T525;
  wire T526;
  wire T527;
  wire T528;
  wire T529;
  wire T530;
  wire T531;
  wire[54:0] T3125;
  wire[30:0] T532;
  wire[30:0] T533;
  wire[8:0] T534;
  wire[4:0] T535;
  wire[3:0] T536;
  wire[21:0] T537;
  wire[4:0] T538;
  wire[16:0] T539;
  wire T540;
  wire T541;
  wire T542;
  wire T543;
  wire flitsAreTail_8;
  wire T544;
  wire T545;
  wire T546;
  wire T547;
  wire[53:0] T548;
  wire T549;
  wire[30:0] T550;
  wire T551;
  wire T552;
  wire T553;
  wire T554;
  wire T555;
  wire[54:0] T556;
  wire[54:0] T557;
  wire T558;
  wire T559;
  wire T560;
  wire T561;
  wire T562;
  wire T563;
  wire T564;
  wire T565;
  wire T566;
  wire T567;
  wire[54:0] T568;
  wire[54:0] T569;
  wire T3126;
  reg [54:0] R570;
  wire[54:0] T3127;
  wire[54:0] T571;
  wire[54:0] T3128;
  wire T572;
  wire T573;
  wire[54:0] T574;
  wire[54:0] T575;
  wire T576;
  wire T577;
  wire[1:0] T578;
  wire[1:0] T579;
  wire[1:0] T580;
  wire T581;
  wire[2:0] T582;
  reg [2:0] R583;
  wire[2:0] T3129;
  wire[1:0] T584;
  wire T585;
  wire T586;
  wire T587;
  wire T588;
  wire T589;
  wire T590;
  wire T591;
  wire T592;
  wire T593;
  wire[2:0] T594;
  wire T595;
  wire T596;
  wire T597;
  wire T598;
  wire T599;
  wire T600;
  wire T601;
  wire T602;
  wire T603;
  wire T604;
  wire T605;
  wire T606;
  wire T607;
  wire T3130;
  wire T608;
  wire T609;
  wire[3:0] T610;
  wire[3:0] T611;
  wire[3:0] T612;
  wire T613;
  wire[2:0] T614;
  wire[3:0] T615;
  wire T616;
  wire T617;
  wire T618;
  wire T619;
  wire T620;
  wire T621;
  wire T622;
  wire[2:0] T623;
  wire T624;
  wire T625;
  wire T626;
  wire T627;
  wire T628;
  wire T629;
  wire T630;
  wire T631;
  wire[53:0] T632;
  wire T633;
  wire[30:0] T634;
  wire T635;
  wire T636;
  reg  R637;
  wire T3131;
  wire[2:0] T638;
  wire[30:0] T639;
  wire[54:0] T640;
  wire[1:0] T641;
  wire[1:0] T642;
  wire[1:0] T643;
  wire[3:0] T644;
  wire T645;
  wire T646;
  wire[15:0] T647;
  wire T648;
  wire T649;
  wire T650;
  wire T651;
  wire T652;
  wire T653;
  wire T654;
  wire T655;
  wire T656;
  wire T657;
  wire T658;
  wire T659;
  wire T660;
  wire T661;
  wire T662;
  wire T663;
  wire T664;
  wire T665;
  wire T666;
  wire T667;
  wire T668;
  wire T669;
  wire T670;
  wire T671;
  wire T672;
  wire T673;
  wire T674;
  wire T675;
  wire[54:0] T3132;
  wire[30:0] T676;
  wire[30:0] T677;
  wire[8:0] T678;
  wire[4:0] T679;
  wire[3:0] T680;
  wire[21:0] T681;
  wire[4:0] T682;
  wire[16:0] T683;
  wire T684;
  wire T685;
  wire T686;
  wire T687;
  wire flitsAreTail_7;
  wire T688;
  wire T689;
  wire T690;
  wire T691;
  wire[53:0] T692;
  wire T693;
  wire[30:0] T694;
  wire T695;
  wire T696;
  wire T697;
  wire T698;
  wire T699;
  wire[54:0] T700;
  wire[54:0] T701;
  wire T702;
  wire T703;
  wire T704;
  wire T705;
  wire T706;
  wire T707;
  wire T708;
  wire T709;
  wire T710;
  wire T711;
  wire[54:0] T712;
  wire[54:0] T713;
  wire T3133;
  reg [54:0] R714;
  wire[54:0] T3134;
  wire[54:0] T715;
  wire[54:0] T3135;
  wire T716;
  wire T717;
  wire[54:0] T718;
  wire[54:0] T719;
  wire T720;
  wire T721;
  wire[1:0] T722;
  wire[1:0] T723;
  wire[1:0] T724;
  wire T725;
  wire[2:0] T726;
  reg [2:0] R727;
  wire[2:0] T3136;
  wire[1:0] T728;
  wire T729;
  wire T730;
  wire T731;
  wire T732;
  wire T733;
  wire T734;
  wire T735;
  wire T736;
  wire T737;
  wire[2:0] T738;
  wire T739;
  wire T740;
  wire T741;
  wire T742;
  wire T743;
  wire T744;
  wire T745;
  wire T746;
  wire T747;
  wire T748;
  wire T749;
  wire T750;
  wire T751;
  wire T3137;
  wire T752;
  wire T753;
  wire[3:0] T754;
  wire[3:0] T755;
  wire[3:0] T756;
  wire T757;
  wire[2:0] T758;
  wire[3:0] T759;
  wire T760;
  wire T761;
  wire T762;
  wire T763;
  wire T764;
  wire T765;
  wire T766;
  wire[2:0] T767;
  wire T768;
  wire T769;
  wire T770;
  wire T771;
  wire T772;
  wire T773;
  wire T774;
  wire T775;
  wire[53:0] T776;
  wire T777;
  wire[30:0] T778;
  wire T779;
  wire T780;
  reg  R781;
  wire T3138;
  wire[2:0] T782;
  wire[30:0] T783;
  wire[54:0] T784;
  wire[1:0] T785;
  wire[1:0] T786;
  wire[1:0] T787;
  wire[3:0] T788;
  wire T789;
  wire T790;
  wire[15:0] T791;
  wire T792;
  wire T793;
  wire T794;
  wire T795;
  wire T796;
  wire T797;
  wire T798;
  wire T799;
  wire T800;
  wire T801;
  wire T802;
  wire T803;
  wire T804;
  wire T805;
  wire T806;
  wire T807;
  wire T808;
  wire T809;
  wire T810;
  wire T811;
  wire T812;
  wire T813;
  wire T814;
  wire T815;
  wire T816;
  wire T817;
  wire T818;
  wire T819;
  wire[54:0] T3139;
  wire[30:0] T820;
  wire[30:0] T821;
  wire[8:0] T822;
  wire[4:0] T823;
  wire[3:0] T824;
  wire[21:0] T825;
  wire[4:0] T826;
  wire[16:0] T827;
  wire T828;
  wire T829;
  wire T830;
  wire T831;
  wire flitsAreTail_6;
  wire T832;
  wire T833;
  wire T834;
  wire T835;
  wire[53:0] T836;
  wire T837;
  wire[30:0] T838;
  wire T839;
  wire T840;
  wire T841;
  wire T842;
  wire T843;
  wire[54:0] T844;
  wire[54:0] T845;
  wire T846;
  wire T847;
  wire T848;
  wire T849;
  wire T850;
  wire T851;
  wire T852;
  wire T853;
  wire T854;
  wire T855;
  wire[54:0] T856;
  wire[54:0] T857;
  wire T3140;
  reg [54:0] R858;
  wire[54:0] T3141;
  wire[54:0] T859;
  wire[54:0] T3142;
  wire T860;
  wire T861;
  wire[54:0] T862;
  wire[54:0] T863;
  wire T864;
  wire T865;
  wire[1:0] T866;
  wire[1:0] T867;
  wire[1:0] T868;
  wire T869;
  wire[2:0] T870;
  reg [2:0] R871;
  wire[2:0] T3143;
  wire[1:0] T872;
  wire T873;
  wire T874;
  wire T875;
  wire T876;
  wire T877;
  wire T878;
  wire T879;
  wire T880;
  wire T881;
  wire[2:0] T882;
  wire T883;
  wire T884;
  wire T885;
  wire T886;
  wire T887;
  wire T888;
  wire T889;
  wire T890;
  wire T891;
  wire T892;
  wire T893;
  wire T894;
  wire T895;
  wire T3144;
  wire T896;
  wire T897;
  wire[3:0] T898;
  wire[3:0] T899;
  wire[3:0] T900;
  wire T901;
  wire[2:0] T902;
  wire[3:0] T903;
  wire T904;
  wire T905;
  wire T906;
  wire T907;
  wire T908;
  wire T909;
  wire T910;
  wire[2:0] T911;
  wire T912;
  wire T913;
  wire T914;
  wire T915;
  wire T916;
  wire T917;
  wire T918;
  wire T919;
  wire[53:0] T920;
  wire T921;
  wire[30:0] T922;
  wire T923;
  wire T924;
  reg  R925;
  wire T3145;
  wire[2:0] T926;
  wire[30:0] T927;
  wire[54:0] T928;
  wire[1:0] T929;
  wire[1:0] T930;
  wire[1:0] T931;
  wire[3:0] T932;
  wire T933;
  wire T934;
  wire[15:0] T935;
  wire T936;
  wire T937;
  wire T938;
  wire T939;
  wire T940;
  wire T941;
  wire T942;
  wire T943;
  wire T944;
  wire T945;
  wire T946;
  wire T947;
  wire T948;
  wire T949;
  wire T950;
  wire T951;
  wire T952;
  wire T953;
  wire T954;
  wire T955;
  wire T956;
  wire T957;
  wire T958;
  wire T959;
  wire T960;
  wire T961;
  wire T962;
  wire T963;
  wire[54:0] T3146;
  wire[30:0] T964;
  wire[30:0] T965;
  wire[8:0] T966;
  wire[4:0] T967;
  wire[3:0] T968;
  wire[21:0] T969;
  wire[4:0] T970;
  wire[16:0] T971;
  wire T972;
  wire T973;
  wire T974;
  wire T975;
  wire flitsAreTail_5;
  wire T976;
  wire T977;
  wire T978;
  wire T979;
  wire[53:0] T980;
  wire T981;
  wire[30:0] T982;
  wire T983;
  wire T984;
  wire T985;
  wire T986;
  wire T987;
  wire[54:0] T988;
  wire[54:0] T989;
  wire T990;
  wire T991;
  wire T992;
  wire T993;
  wire T994;
  wire T995;
  wire T996;
  wire T997;
  wire T998;
  wire T999;
  wire[54:0] T1000;
  wire[54:0] T1001;
  wire T3147;
  reg [54:0] R1002;
  wire[54:0] T3148;
  wire[54:0] T1003;
  wire[54:0] T3149;
  wire T1004;
  wire T1005;
  wire[54:0] T1006;
  wire[54:0] T1007;
  wire T1008;
  wire T1009;
  wire[1:0] T1010;
  wire[1:0] T1011;
  wire[1:0] T1012;
  wire T1013;
  wire[2:0] T1014;
  reg [2:0] R1015;
  wire[2:0] T3150;
  wire[1:0] T1016;
  wire T1017;
  wire T1018;
  wire T1019;
  wire T1020;
  wire T1021;
  wire T1022;
  wire T1023;
  wire T1024;
  wire T1025;
  wire[2:0] T1026;
  wire T1027;
  wire T1028;
  wire T1029;
  wire T1030;
  wire T1031;
  wire T1032;
  wire T1033;
  wire T1034;
  wire T1035;
  wire T1036;
  wire T1037;
  wire T1038;
  wire T1039;
  wire T3151;
  wire T1040;
  wire T1041;
  wire[3:0] T1042;
  wire[3:0] T1043;
  wire[3:0] T1044;
  wire T1045;
  wire[2:0] T1046;
  wire[3:0] T1047;
  wire T1048;
  wire T1049;
  wire T1050;
  wire T1051;
  wire T1052;
  wire T1053;
  wire T1054;
  wire[2:0] T1055;
  wire T1056;
  wire T1057;
  wire T1058;
  wire T1059;
  wire T1060;
  wire T1061;
  wire T1062;
  wire T1063;
  wire[53:0] T1064;
  wire T1065;
  wire[30:0] T1066;
  wire T1067;
  wire T1068;
  reg  R1069;
  wire T3152;
  wire[2:0] T1070;
  wire[30:0] T1071;
  wire[54:0] T1072;
  wire[1:0] T1073;
  wire[1:0] T1074;
  wire[1:0] T1075;
  wire[3:0] T1076;
  wire T1077;
  wire T1078;
  wire[15:0] T1079;
  wire T1080;
  wire T1081;
  wire T1082;
  wire T1083;
  wire T1084;
  wire T1085;
  wire T1086;
  wire T1087;
  wire T1088;
  wire T1089;
  wire T1090;
  wire T1091;
  wire T1092;
  wire T1093;
  wire T1094;
  wire T1095;
  wire T1096;
  wire T1097;
  wire T1098;
  wire T1099;
  wire T1100;
  wire T1101;
  wire T1102;
  wire T1103;
  wire T1104;
  wire T1105;
  wire T1106;
  wire T1107;
  wire[54:0] T3153;
  wire[30:0] T1108;
  wire[30:0] T1109;
  wire[8:0] T1110;
  wire[4:0] T1111;
  wire[3:0] T1112;
  wire[21:0] T1113;
  wire[4:0] T1114;
  wire[16:0] T1115;
  wire T1116;
  wire T1117;
  wire T1118;
  wire T1119;
  wire flitsAreTail_4;
  wire T1120;
  wire T1121;
  wire T1122;
  wire T1123;
  wire[53:0] T1124;
  wire T1125;
  wire[30:0] T1126;
  wire T1127;
  wire T1128;
  wire T1129;
  wire T1130;
  wire T1131;
  wire[54:0] T1132;
  wire[54:0] T1133;
  wire T1134;
  wire T1135;
  wire T1136;
  wire T1137;
  wire T1138;
  wire T1139;
  wire T1140;
  wire T1141;
  wire T1142;
  wire T1143;
  wire[54:0] T1144;
  wire[54:0] T1145;
  wire T3154;
  reg [54:0] R1146;
  wire[54:0] T3155;
  wire[54:0] T1147;
  wire[54:0] T3156;
  wire T1148;
  wire T1149;
  wire[54:0] T1150;
  wire[54:0] T1151;
  wire T1152;
  wire T1153;
  wire[1:0] T1154;
  wire[1:0] T1155;
  wire[1:0] T1156;
  wire T1157;
  wire[2:0] T1158;
  reg [2:0] R1159;
  wire[2:0] T3157;
  wire[1:0] T1160;
  wire T1161;
  wire T1162;
  wire T1163;
  wire T1164;
  wire T1165;
  wire T1166;
  wire T1167;
  wire T1168;
  wire T1169;
  wire[2:0] T1170;
  wire T1171;
  wire T1172;
  wire T1173;
  wire T1174;
  wire T1175;
  wire T1176;
  wire T1177;
  wire T1178;
  wire T1179;
  wire T1180;
  wire T1181;
  wire T1182;
  wire T1183;
  wire T3158;
  wire T1184;
  wire T1185;
  wire[3:0] T1186;
  wire[3:0] T1187;
  wire[3:0] T1188;
  wire T1189;
  wire[2:0] T1190;
  wire[3:0] T1191;
  wire T1192;
  wire T1193;
  wire T1194;
  wire T1195;
  wire T1196;
  wire T1197;
  wire T1198;
  wire[2:0] T1199;
  wire T1200;
  wire T1201;
  wire T1202;
  wire T1203;
  wire T1204;
  wire T1205;
  wire T1206;
  wire T1207;
  wire[53:0] T1208;
  wire T1209;
  wire[30:0] T1210;
  wire T1211;
  wire T1212;
  reg  R1213;
  wire T3159;
  wire[2:0] T1214;
  wire[30:0] T1215;
  wire[54:0] T1216;
  wire[1:0] T1217;
  wire[1:0] T1218;
  wire[1:0] T1219;
  wire[3:0] T1220;
  wire T1221;
  wire T1222;
  wire[15:0] T1223;
  wire T1224;
  wire T1225;
  wire T1226;
  wire T1227;
  wire T1228;
  wire T1229;
  wire T1230;
  wire T1231;
  wire T1232;
  wire T1233;
  wire T1234;
  wire T1235;
  wire T1236;
  wire T1237;
  wire T1238;
  wire T1239;
  wire T1240;
  wire T1241;
  wire T1242;
  wire T1243;
  wire T1244;
  wire T1245;
  wire T1246;
  wire T1247;
  wire T1248;
  wire T1249;
  wire T1250;
  wire T1251;
  wire[54:0] T3160;
  wire[30:0] T1252;
  wire[30:0] T1253;
  wire[8:0] T1254;
  wire[4:0] T1255;
  wire[3:0] T1256;
  wire[21:0] T1257;
  wire[4:0] T1258;
  wire[16:0] T1259;
  wire T1260;
  wire T1261;
  wire T1262;
  wire T1263;
  wire flitsAreTail_3;
  wire T1264;
  wire T1265;
  wire T1266;
  wire T1267;
  wire[53:0] T1268;
  wire T1269;
  wire[30:0] T1270;
  wire T1271;
  wire T1272;
  wire T1273;
  wire T1274;
  wire T1275;
  wire[54:0] T1276;
  wire[54:0] T1277;
  wire T1278;
  wire T1279;
  wire T1280;
  wire T1281;
  wire T1282;
  wire T1283;
  wire T1284;
  wire T1285;
  wire T1286;
  wire T1287;
  wire[54:0] T1288;
  wire[54:0] T1289;
  wire T3161;
  reg [54:0] R1290;
  wire[54:0] T3162;
  wire[54:0] T1291;
  wire[54:0] T3163;
  wire T1292;
  wire T1293;
  wire[54:0] T1294;
  wire[54:0] T1295;
  wire T1296;
  wire T1297;
  wire[1:0] T1298;
  wire[1:0] T1299;
  wire[1:0] T1300;
  wire T1301;
  wire[2:0] T1302;
  reg [2:0] R1303;
  wire[2:0] T3164;
  wire[1:0] T1304;
  wire T1305;
  wire T1306;
  wire T1307;
  wire T1308;
  wire T1309;
  wire T1310;
  wire T1311;
  wire T1312;
  wire T1313;
  wire[2:0] T1314;
  wire T1315;
  wire T1316;
  wire T1317;
  wire T1318;
  wire T1319;
  wire T1320;
  wire T1321;
  wire T1322;
  wire T1323;
  wire T1324;
  wire T1325;
  wire T1326;
  wire T1327;
  wire T3165;
  wire T1328;
  wire T1329;
  wire[3:0] T1330;
  wire[3:0] T1331;
  wire[3:0] T1332;
  wire T1333;
  wire[2:0] T1334;
  wire[3:0] T1335;
  wire T1336;
  wire T1337;
  wire T1338;
  wire T1339;
  wire T1340;
  wire T1341;
  wire T1342;
  wire[2:0] T1343;
  wire T1344;
  wire T1345;
  wire T1346;
  wire T1347;
  wire T1348;
  wire T1349;
  wire T1350;
  wire T1351;
  wire[53:0] T1352;
  wire T1353;
  wire[30:0] T1354;
  wire T1355;
  wire T1356;
  reg  R1357;
  wire T3166;
  wire[2:0] T1358;
  wire[30:0] T1359;
  wire[54:0] T1360;
  wire[1:0] T1361;
  wire[1:0] T1362;
  wire[1:0] T1363;
  wire[3:0] T1364;
  wire T1365;
  wire T1366;
  wire[15:0] T1367;
  wire T1368;
  wire T1369;
  wire T1370;
  wire T1371;
  wire T1372;
  wire T1373;
  wire T1374;
  wire T1375;
  wire T1376;
  wire T1377;
  wire T1378;
  wire T1379;
  wire T1380;
  wire T1381;
  wire T1382;
  wire T1383;
  wire T1384;
  wire T1385;
  wire T1386;
  wire T1387;
  wire T1388;
  wire T1389;
  wire T1390;
  wire T1391;
  wire T1392;
  wire T1393;
  wire T1394;
  wire T1395;
  wire[54:0] T3167;
  wire[30:0] T1396;
  wire[30:0] T1397;
  wire[8:0] T1398;
  wire[4:0] T1399;
  wire[3:0] T1400;
  wire[21:0] T1401;
  wire[4:0] T1402;
  wire[16:0] T1403;
  wire T1404;
  wire T1405;
  wire T1406;
  wire T1407;
  wire flitsAreTail_2;
  wire T1408;
  wire T1409;
  wire T1410;
  wire T1411;
  wire[53:0] T1412;
  wire T1413;
  wire[30:0] T1414;
  wire T1415;
  wire T1416;
  wire T1417;
  wire T1418;
  wire T1419;
  wire[54:0] T1420;
  wire[54:0] T1421;
  wire T1422;
  wire T1423;
  wire T1424;
  wire T1425;
  wire T1426;
  wire T1427;
  wire T1428;
  wire T1429;
  wire T1430;
  wire T1431;
  wire[54:0] T1432;
  wire[54:0] T1433;
  wire T3168;
  reg [54:0] R1434;
  wire[54:0] T3169;
  wire[54:0] T1435;
  wire[54:0] T3170;
  wire T1436;
  wire T1437;
  wire[54:0] T1438;
  wire[54:0] T1439;
  wire T1440;
  wire T1441;
  wire[1:0] T1442;
  wire[1:0] T1443;
  wire[1:0] T1444;
  wire T1445;
  wire[2:0] T1446;
  reg [2:0] R1447;
  wire[2:0] T3171;
  wire[1:0] T1448;
  wire T1449;
  wire T1450;
  wire T1451;
  wire T1452;
  wire T1453;
  wire T1454;
  wire T1455;
  wire T1456;
  wire T1457;
  wire[2:0] T1458;
  wire T1459;
  wire T1460;
  wire T1461;
  wire T1462;
  wire T1463;
  wire T1464;
  wire T1465;
  wire T1466;
  wire T1467;
  wire T1468;
  wire T1469;
  wire T1470;
  wire T1471;
  wire T3172;
  wire T1472;
  wire T1473;
  wire[3:0] T1474;
  wire[3:0] T1475;
  wire[3:0] T1476;
  wire T1477;
  wire[2:0] T1478;
  wire[3:0] T1479;
  wire T1480;
  wire T1481;
  wire T1482;
  wire T1483;
  wire T1484;
  wire T1485;
  wire T1486;
  wire[2:0] T1487;
  wire T1488;
  wire T1489;
  wire T1490;
  wire T1491;
  wire T1492;
  wire T1493;
  wire T1494;
  wire T1495;
  wire[53:0] T1496;
  wire T1497;
  wire[30:0] T1498;
  wire T1499;
  wire T1500;
  reg  R1501;
  wire T3173;
  wire[2:0] T1502;
  wire[30:0] T1503;
  wire[54:0] T1504;
  wire[1:0] T1505;
  wire[1:0] T1506;
  wire[1:0] T1507;
  wire[3:0] T1508;
  wire T1509;
  wire T1510;
  wire[15:0] T1511;
  wire T1512;
  wire T1513;
  wire T1514;
  wire T1515;
  wire T1516;
  wire T1517;
  wire T1518;
  wire T1519;
  wire T1520;
  wire T1521;
  wire T1522;
  wire T1523;
  wire T1524;
  wire T1525;
  wire T1526;
  wire T1527;
  wire T1528;
  wire T1529;
  wire T1530;
  wire T1531;
  wire T1532;
  wire T1533;
  wire T1534;
  wire T1535;
  wire T1536;
  wire T1537;
  wire T1538;
  wire T1539;
  wire[54:0] T3174;
  wire[30:0] T1540;
  wire[30:0] T1541;
  wire[8:0] T1542;
  wire[4:0] T1543;
  wire[3:0] T1544;
  wire[21:0] T1545;
  wire[4:0] T1546;
  wire[16:0] T1547;
  wire T1548;
  wire T1549;
  wire T1550;
  wire T1551;
  wire flitsAreTail_1;
  wire T1552;
  wire T1553;
  wire T1554;
  wire T1555;
  wire[53:0] T1556;
  wire T1557;
  wire[30:0] T1558;
  wire T1559;
  wire T1560;
  wire T1561;
  wire T1562;
  wire T1563;
  wire[54:0] T1564;
  wire[54:0] T1565;
  wire T1566;
  wire T1567;
  wire T1568;
  wire T1569;
  wire T1570;
  wire T1571;
  wire T1572;
  wire T1573;
  wire T1574;
  wire T1575;
  wire[54:0] T1576;
  wire[54:0] T1577;
  wire T3175;
  reg [54:0] R1578;
  wire[54:0] T3176;
  wire[54:0] T1579;
  wire[54:0] T3177;
  wire T1580;
  wire T1581;
  wire[54:0] T1582;
  wire[54:0] T1583;
  wire T1584;
  wire T1585;
  wire[1:0] T1586;
  wire[1:0] T1587;
  wire[1:0] T1588;
  wire T1589;
  wire[2:0] T1590;
  reg [2:0] R1591;
  wire[2:0] T3178;
  wire[1:0] T1592;
  wire T1593;
  wire T1594;
  wire T1595;
  wire T1596;
  wire T1597;
  wire T1598;
  wire T1599;
  wire T1600;
  wire T1601;
  wire[2:0] T1602;
  wire T1603;
  wire T1604;
  wire T1605;
  wire T1606;
  wire T1607;
  wire T1608;
  wire T1609;
  wire T1610;
  wire T1611;
  wire T1612;
  wire T1613;
  wire T1614;
  wire T1615;
  wire T3179;
  wire T1616;
  wire T1617;
  wire[3:0] T1618;
  wire[3:0] T1619;
  wire[3:0] T1620;
  wire T1621;
  wire[2:0] T1622;
  wire[3:0] T1623;
  wire T1624;
  wire T1625;
  wire T1626;
  wire T1627;
  wire T1628;
  wire T1629;
  wire T1630;
  wire[2:0] T1631;
  wire T1632;
  wire T1633;
  wire T1634;
  wire T1635;
  wire T1636;
  wire T1637;
  wire T1638;
  wire T1639;
  wire[53:0] T1640;
  wire T1641;
  wire[30:0] T1642;
  wire T1643;
  wire T1644;
  reg  R1645;
  wire T3180;
  wire[2:0] T1646;
  wire[30:0] T1647;
  wire[54:0] T1648;
  wire[1:0] T1649;
  wire[1:0] T1650;
  wire[1:0] T1651;
  wire[3:0] T1652;
  wire T1653;
  wire T1654;
  wire[15:0] T1655;
  wire T1656;
  wire T1657;
  wire T1658;
  wire T1659;
  wire T1660;
  wire T1661;
  wire T1662;
  wire T1663;
  wire T1664;
  wire T1665;
  wire T1666;
  wire T1667;
  wire T1668;
  wire T1669;
  wire T1670;
  wire T1671;
  wire T1672;
  wire T1673;
  wire T1674;
  wire T1675;
  wire T1676;
  wire T1677;
  wire T1678;
  wire T1679;
  wire T1680;
  wire T1681;
  wire T1682;
  wire T1683;
  wire[54:0] T3181;
  wire[30:0] T1684;
  wire[30:0] T1685;
  wire[8:0] T1686;
  wire[4:0] T1687;
  wire[3:0] T1688;
  wire[21:0] T1689;
  wire[4:0] T1690;
  wire[16:0] T1691;
  wire T1692;
  wire T1693;
  wire T1694;
  wire T1695;
  wire flitsAreTail_0;
  wire T1696;
  wire T1697;
  wire T1698;
  wire T1699;
  wire[53:0] T1700;
  wire T1701;
  wire[30:0] T1702;
  wire T1703;
  wire T1704;
  wire T1705;
  wire T1706;
  wire T1707;
  wire[54:0] T1708;
  wire[54:0] T1709;
  wire T1710;
  wire T1711;
  wire T1712;
  wire T1713;
  wire T1714;
  wire T1715;
  wire T1716;
  wire T1717;
  wire T1718;
  wire T1719;
  wire T1720;
  wire T1721;
  wire T1722;
  wire[9:0] T1723;
  wire[9:0] T1724;
  wire[4:0] T1725;
  wire[2:0] T1726;
  wire[1:0] T1727;
  wire readyToXmit_0_4;
  wire T1728;
  wire T1729;
  wire T1730;
  wire T1731;
  wire T1732;
  wire T1733;
  wire T1734;
  wire T1735;
  wire[7:0] T1736;
  wire[2:0] T1737;
  wire T1738;
  wire T1739;
  wire T1740;
  wire T1741;
  wire T1742;
  wire T1743;
  wire T1744;
  wire readyToXmit_1_4;
  wire T1745;
  wire T1746;
  wire T1747;
  wire T1748;
  wire T1749;
  wire T1750;
  wire T1751;
  wire T1752;
  wire[7:0] T1753;
  wire[2:0] T1754;
  wire T1755;
  wire T1756;
  wire T1757;
  wire T1758;
  wire T1759;
  wire T1760;
  wire T1761;
  wire readyToXmit_2_4;
  wire T1762;
  wire T1763;
  wire T1764;
  wire T1765;
  wire T1766;
  wire T1767;
  wire T1768;
  wire T1769;
  wire[7:0] T1770;
  wire[2:0] T1771;
  wire T1772;
  wire T1773;
  wire T1774;
  wire T1775;
  wire T1776;
  wire T1777;
  wire T1778;
  wire[1:0] T1779;
  wire readyToXmit_3_4;
  wire T1780;
  wire T1781;
  wire T1782;
  wire T1783;
  wire T1784;
  wire T1785;
  wire T1786;
  wire T1787;
  wire[7:0] T1788;
  wire[2:0] T1789;
  wire T1790;
  wire T1791;
  wire T1792;
  wire T1793;
  wire T1794;
  wire T1795;
  wire T1796;
  wire readyToXmit_4_4;
  wire T1797;
  wire T1798;
  wire T1799;
  wire T1800;
  wire T1801;
  wire T1802;
  wire T1803;
  wire T1804;
  wire[7:0] T1805;
  wire[2:0] T1806;
  wire T1807;
  wire T1808;
  wire T1809;
  wire T1810;
  wire T1811;
  wire T1812;
  wire T1813;
  wire[4:0] T1814;
  wire[2:0] T1815;
  wire[1:0] T1816;
  wire readyToXmit_5_4;
  wire T1817;
  wire T1818;
  wire T1819;
  wire T1820;
  wire T1821;
  wire T1822;
  wire T1823;
  wire T1824;
  wire[7:0] T1825;
  wire[2:0] T1826;
  wire T1827;
  wire T1828;
  wire T1829;
  wire T1830;
  wire T1831;
  wire T1832;
  wire T1833;
  wire readyToXmit_6_4;
  wire T1834;
  wire T1835;
  wire T1836;
  wire T1837;
  wire T1838;
  wire T1839;
  wire T1840;
  wire T1841;
  wire[7:0] T1842;
  wire[2:0] T1843;
  wire T1844;
  wire T1845;
  wire T1846;
  wire T1847;
  wire T1848;
  wire T1849;
  wire T1850;
  wire readyToXmit_7_4;
  wire T1851;
  wire T1852;
  wire T1853;
  wire T1854;
  wire T1855;
  wire T1856;
  wire T1857;
  wire T1858;
  wire[7:0] T1859;
  wire[2:0] T1860;
  wire T1861;
  wire T1862;
  wire T1863;
  wire T1864;
  wire T1865;
  wire T1866;
  wire T1867;
  wire[1:0] T1868;
  wire readyToXmit_8_4;
  wire T1869;
  wire T1870;
  wire T1871;
  wire T1872;
  wire T1873;
  wire T1874;
  wire T1875;
  wire T1876;
  wire[7:0] T1877;
  wire[2:0] T1878;
  wire T1879;
  wire T1880;
  wire T1881;
  wire T1882;
  wire T1883;
  wire T1884;
  wire T1885;
  wire readyToXmit_9_4;
  wire T1886;
  wire T1887;
  wire T1888;
  wire T1889;
  wire T1890;
  wire T1891;
  wire T1892;
  wire T1893;
  wire[7:0] T1894;
  wire[2:0] T1895;
  wire T1896;
  wire T1897;
  wire T1898;
  wire T1899;
  wire T1900;
  wire T1901;
  wire T1902;
  wire T1903;
  wire T1904;
  wire T1905;
  wire[9:0] T1906;
  wire[9:0] T1907;
  wire[4:0] T1908;
  wire[2:0] T1909;
  wire[1:0] T1910;
  wire readyToXmit_0_3;
  wire T1911;
  wire T1912;
  wire T1913;
  wire T1914;
  wire T1915;
  wire readyToXmit_1_3;
  wire T1916;
  wire T1917;
  wire T1918;
  wire T1919;
  wire T1920;
  wire readyToXmit_2_3;
  wire T1921;
  wire T1922;
  wire T1923;
  wire T1924;
  wire T1925;
  wire[1:0] T1926;
  wire readyToXmit_3_3;
  wire T1927;
  wire T1928;
  wire T1929;
  wire T1930;
  wire T1931;
  wire readyToXmit_4_3;
  wire T1932;
  wire T1933;
  wire T1934;
  wire T1935;
  wire T1936;
  wire[4:0] T1937;
  wire[2:0] T1938;
  wire[1:0] T1939;
  wire readyToXmit_5_3;
  wire T1940;
  wire T1941;
  wire T1942;
  wire T1943;
  wire T1944;
  wire readyToXmit_6_3;
  wire T1945;
  wire T1946;
  wire T1947;
  wire T1948;
  wire T1949;
  wire readyToXmit_7_3;
  wire T1950;
  wire T1951;
  wire T1952;
  wire T1953;
  wire T1954;
  wire[1:0] T1955;
  wire readyToXmit_8_3;
  wire T1956;
  wire T1957;
  wire T1958;
  wire T1959;
  wire T1960;
  wire readyToXmit_9_3;
  wire T1961;
  wire T1962;
  wire T1963;
  wire T1964;
  wire T1965;
  wire T1966;
  wire T1967;
  wire T1968;
  wire[9:0] T1969;
  wire[9:0] T1970;
  wire[4:0] T1971;
  wire[2:0] T1972;
  wire[1:0] T1973;
  wire readyToXmit_0_2;
  wire T1974;
  wire T1975;
  wire T1976;
  wire T1977;
  wire T1978;
  wire readyToXmit_1_2;
  wire T1979;
  wire T1980;
  wire T1981;
  wire T1982;
  wire T1983;
  wire readyToXmit_2_2;
  wire T1984;
  wire T1985;
  wire T1986;
  wire T1987;
  wire T1988;
  wire[1:0] T1989;
  wire readyToXmit_3_2;
  wire T1990;
  wire T1991;
  wire T1992;
  wire T1993;
  wire T1994;
  wire readyToXmit_4_2;
  wire T1995;
  wire T1996;
  wire T1997;
  wire T1998;
  wire T1999;
  wire[4:0] T2000;
  wire[2:0] T2001;
  wire[1:0] T2002;
  wire readyToXmit_5_2;
  wire T2003;
  wire T2004;
  wire T2005;
  wire T2006;
  wire T2007;
  wire readyToXmit_6_2;
  wire T2008;
  wire T2009;
  wire T2010;
  wire T2011;
  wire T2012;
  wire readyToXmit_7_2;
  wire T2013;
  wire T2014;
  wire T2015;
  wire T2016;
  wire T2017;
  wire[1:0] T2018;
  wire readyToXmit_8_2;
  wire T2019;
  wire T2020;
  wire T2021;
  wire T2022;
  wire T2023;
  wire readyToXmit_9_2;
  wire T2024;
  wire T2025;
  wire T2026;
  wire T2027;
  wire T2028;
  wire T2029;
  wire T2030;
  wire T2031;
  wire[9:0] T2032;
  wire[9:0] T2033;
  wire[4:0] T2034;
  wire[2:0] T2035;
  wire[1:0] T2036;
  wire readyToXmit_0_1;
  wire T2037;
  wire T2038;
  wire T2039;
  wire T2040;
  wire T2041;
  wire readyToXmit_1_1;
  wire T2042;
  wire T2043;
  wire T2044;
  wire T2045;
  wire T2046;
  wire readyToXmit_2_1;
  wire T2047;
  wire T2048;
  wire T2049;
  wire T2050;
  wire T2051;
  wire[1:0] T2052;
  wire readyToXmit_3_1;
  wire T2053;
  wire T2054;
  wire T2055;
  wire T2056;
  wire T2057;
  wire readyToXmit_4_1;
  wire T2058;
  wire T2059;
  wire T2060;
  wire T2061;
  wire T2062;
  wire[4:0] T2063;
  wire[2:0] T2064;
  wire[1:0] T2065;
  wire readyToXmit_5_1;
  wire T2066;
  wire T2067;
  wire T2068;
  wire T2069;
  wire T2070;
  wire readyToXmit_6_1;
  wire T2071;
  wire T2072;
  wire T2073;
  wire T2074;
  wire T2075;
  wire readyToXmit_7_1;
  wire T2076;
  wire T2077;
  wire T2078;
  wire T2079;
  wire T2080;
  wire[1:0] T2081;
  wire readyToXmit_8_1;
  wire T2082;
  wire T2083;
  wire T2084;
  wire T2085;
  wire T2086;
  wire readyToXmit_9_1;
  wire T2087;
  wire T2088;
  wire T2089;
  wire T2090;
  wire T2091;
  wire T2092;
  wire T2093;
  wire T2094;
  wire[9:0] T2095;
  wire[9:0] T2096;
  wire[4:0] T2097;
  wire[2:0] T2098;
  wire[1:0] T2099;
  wire readyToXmit_0_0;
  wire T2100;
  wire T2101;
  wire T2102;
  wire T2103;
  wire T2104;
  wire readyToXmit_1_0;
  wire T2105;
  wire T2106;
  wire T2107;
  wire T2108;
  wire T2109;
  wire readyToXmit_2_0;
  wire T2110;
  wire T2111;
  wire T2112;
  wire T2113;
  wire T2114;
  wire[1:0] T2115;
  wire readyToXmit_3_0;
  wire T2116;
  wire T2117;
  wire T2118;
  wire T2119;
  wire T2120;
  wire readyToXmit_4_0;
  wire T2121;
  wire T2122;
  wire T2123;
  wire T2124;
  wire T2125;
  wire[4:0] T2126;
  wire[2:0] T2127;
  wire[1:0] T2128;
  wire readyToXmit_5_0;
  wire T2129;
  wire T2130;
  wire T2131;
  wire T2132;
  wire T2133;
  wire readyToXmit_6_0;
  wire T2134;
  wire T2135;
  wire T2136;
  wire T2137;
  wire T2138;
  wire readyToXmit_7_0;
  wire T2139;
  wire T2140;
  wire T2141;
  wire T2142;
  wire T2143;
  wire[1:0] T2144;
  wire readyToXmit_8_0;
  wire T2145;
  wire T2146;
  wire T2147;
  wire T2148;
  wire T2149;
  wire readyToXmit_9_0;
  wire T2150;
  wire T2151;
  wire T2152;
  wire T2153;
  wire T2154;
  wire T2155;
  wire T2156;
  wire T2157;
  wire T2158;
  wire T2159;
  wire T2160;
  wire T2161;
  wire T2162;
  wire T2163;
  wire T2164;
  wire T2165;
  wire T2166;
  wire T2167;
  wire T2168;
  wire T2169;
  wire T2170;
  wire T2171;
  wire T2172;
  wire T2173;
  wire T2174;
  wire T2175;
  reg [1:0] validVCs_0_0;
  reg  R2176;
  wire T2177;
  wire T2178;
  wire T2179;
  wire T2180;
  reg  R2181;
  wire T2182;
  wire T2183;
  wire T2184;
  wire T2185;
  reg [1:0] validVCs_0_1;
  reg  R2186;
  wire T2187;
  wire T2188;
  wire T2189;
  wire T2190;
  reg  R2191;
  wire T2192;
  wire T2193;
  wire T2194;
  wire T2195;
  reg [1:0] validVCs_0_2;
  reg  R2196;
  wire T2197;
  wire T2198;
  wire T2199;
  wire T2200;
  reg  R2201;
  wire T2202;
  wire T2203;
  wire T2204;
  wire T2205;
  reg [1:0] validVCs_0_3;
  reg  R2206;
  wire T2207;
  wire T2208;
  wire T2209;
  wire T2210;
  reg  R2211;
  wire T2212;
  wire T2213;
  wire T2214;
  wire T2215;
  reg [1:0] validVCs_0_4;
  reg  R2216;
  wire T2217;
  wire T2218;
  wire T2219;
  wire T2220;
  reg  R2221;
  wire T2222;
  wire T2223;
  wire T2224;
  wire T2225;
  reg [1:0] validVCs_1_0;
  reg  R2226;
  wire T2227;
  wire T2228;
  wire T2229;
  wire T2230;
  reg  R2231;
  wire T2232;
  wire T2233;
  wire T2234;
  wire T2235;
  reg [1:0] validVCs_1_1;
  reg  R2236;
  wire T2237;
  wire T2238;
  wire T2239;
  wire T2240;
  reg  R2241;
  wire T2242;
  wire T2243;
  wire T2244;
  wire T2245;
  reg [1:0] validVCs_1_2;
  reg  R2246;
  wire T2247;
  wire T2248;
  wire T2249;
  wire T2250;
  reg  R2251;
  wire T2252;
  wire T2253;
  wire T2254;
  wire T2255;
  reg [1:0] validVCs_1_3;
  reg  R2256;
  wire T2257;
  wire T2258;
  wire T2259;
  wire T2260;
  reg  R2261;
  wire T2262;
  wire T2263;
  wire T2264;
  wire T2265;
  reg [1:0] validVCs_1_4;
  reg  R2266;
  wire T2267;
  wire T2268;
  wire T2269;
  wire T2270;
  reg  R2271;
  wire T2272;
  wire T2273;
  wire T2274;
  wire T2275;
  reg [1:0] validVCs_2_0;
  reg  R2276;
  wire T2277;
  wire T2278;
  wire T2279;
  wire T2280;
  reg  R2281;
  wire T2282;
  wire T2283;
  wire T2284;
  wire T2285;
  reg [1:0] validVCs_2_1;
  reg  R2286;
  wire T2287;
  wire T2288;
  wire T2289;
  wire T2290;
  reg  R2291;
  wire T2292;
  wire T2293;
  wire T2294;
  wire T2295;
  reg [1:0] validVCs_2_2;
  reg  R2296;
  wire T2297;
  wire T2298;
  wire T2299;
  wire T2300;
  reg  R2301;
  wire T2302;
  wire T2303;
  wire T2304;
  wire T2305;
  reg [1:0] validVCs_2_3;
  reg  R2306;
  wire T2307;
  wire T2308;
  wire T2309;
  wire T2310;
  reg  R2311;
  wire T2312;
  wire T2313;
  wire T2314;
  wire T2315;
  reg [1:0] validVCs_2_4;
  reg  R2316;
  wire T2317;
  wire T2318;
  wire T2319;
  wire T2320;
  reg  R2321;
  wire T2322;
  wire T2323;
  wire T2324;
  wire T2325;
  reg [1:0] validVCs_3_0;
  reg  R2326;
  wire T2327;
  wire T2328;
  wire T2329;
  wire T2330;
  reg  R2331;
  wire T2332;
  wire T2333;
  wire T2334;
  wire T2335;
  reg [1:0] validVCs_3_1;
  reg  R2336;
  wire T2337;
  wire T2338;
  wire T2339;
  wire T2340;
  reg  R2341;
  wire T2342;
  wire T2343;
  wire T2344;
  wire T2345;
  reg [1:0] validVCs_3_2;
  reg  R2346;
  wire T2347;
  wire T2348;
  wire T2349;
  wire T2350;
  reg  R2351;
  wire T2352;
  wire T2353;
  wire T2354;
  wire T2355;
  reg [1:0] validVCs_3_3;
  reg  R2356;
  wire T2357;
  wire T2358;
  wire T2359;
  wire T2360;
  reg  R2361;
  wire T2362;
  wire T2363;
  wire T2364;
  wire T2365;
  reg [1:0] validVCs_3_4;
  reg  R2366;
  wire T2367;
  wire T2368;
  wire T2369;
  wire T2370;
  reg  R2371;
  wire T2372;
  wire T2373;
  wire T2374;
  wire T2375;
  reg [1:0] validVCs_4_0;
  reg  R2376;
  wire T2377;
  wire T2378;
  wire T2379;
  wire T2380;
  reg  R2381;
  wire T2382;
  wire T2383;
  wire T2384;
  wire T2385;
  reg [1:0] validVCs_4_1;
  reg  R2386;
  wire T2387;
  wire T2388;
  wire T2389;
  wire T2390;
  reg  R2391;
  wire T2392;
  wire T2393;
  wire T2394;
  wire T2395;
  reg [1:0] validVCs_4_2;
  reg  R2396;
  wire T2397;
  wire T2398;
  wire T2399;
  wire T2400;
  reg  R2401;
  wire T2402;
  wire T2403;
  wire T2404;
  wire T2405;
  reg [1:0] validVCs_4_3;
  reg  R2406;
  wire T2407;
  wire T2408;
  wire T2409;
  wire T2410;
  reg  R2411;
  wire T2412;
  wire T2413;
  wire T2414;
  wire T2415;
  reg [1:0] validVCs_4_4;
  reg  R2416;
  wire T2417;
  wire T2418;
  wire T2419;
  wire T2420;
  reg  R2421;
  wire T2422;
  wire T2423;
  wire T2424;
  wire T2425;
  reg [1:0] validVCs_5_0;
  reg  R2426;
  wire T2427;
  wire T2428;
  wire T2429;
  wire T2430;
  reg  R2431;
  wire T2432;
  wire T2433;
  wire T2434;
  wire T2435;
  reg [1:0] validVCs_5_1;
  reg  R2436;
  wire T2437;
  wire T2438;
  wire T2439;
  wire T2440;
  reg  R2441;
  wire T2442;
  wire T2443;
  wire T2444;
  wire T2445;
  reg [1:0] validVCs_5_2;
  reg  R2446;
  wire T2447;
  wire T2448;
  wire T2449;
  wire T2450;
  reg  R2451;
  wire T2452;
  wire T2453;
  wire T2454;
  wire T2455;
  reg [1:0] validVCs_5_3;
  reg  R2456;
  wire T2457;
  wire T2458;
  wire T2459;
  wire T2460;
  reg  R2461;
  wire T2462;
  wire T2463;
  wire T2464;
  wire T2465;
  reg [1:0] validVCs_5_4;
  reg  R2466;
  wire T2467;
  wire T2468;
  wire T2469;
  wire T2470;
  reg  R2471;
  wire T2472;
  wire T2473;
  wire T2474;
  wire T2475;
  reg [1:0] validVCs_6_0;
  reg  R2476;
  wire T2477;
  wire T2478;
  wire T2479;
  wire T2480;
  reg  R2481;
  wire T2482;
  wire T2483;
  wire T2484;
  wire T2485;
  reg [1:0] validVCs_6_1;
  reg  R2486;
  wire T2487;
  wire T2488;
  wire T2489;
  wire T2490;
  reg  R2491;
  wire T2492;
  wire T2493;
  wire T2494;
  wire T2495;
  reg [1:0] validVCs_6_2;
  reg  R2496;
  wire T2497;
  wire T2498;
  wire T2499;
  wire T2500;
  reg  R2501;
  wire T2502;
  wire T2503;
  wire T2504;
  wire T2505;
  reg [1:0] validVCs_6_3;
  reg  R2506;
  wire T2507;
  wire T2508;
  wire T2509;
  wire T2510;
  reg  R2511;
  wire T2512;
  wire T2513;
  wire T2514;
  wire T2515;
  reg [1:0] validVCs_6_4;
  reg  R2516;
  wire T2517;
  wire T2518;
  wire T2519;
  wire T2520;
  reg  R2521;
  wire T2522;
  wire T2523;
  wire T2524;
  wire T2525;
  reg [1:0] validVCs_7_0;
  reg  R2526;
  wire T2527;
  wire T2528;
  wire T2529;
  wire T2530;
  reg  R2531;
  wire T2532;
  wire T2533;
  wire T2534;
  wire T2535;
  reg [1:0] validVCs_7_1;
  reg  R2536;
  wire T2537;
  wire T2538;
  wire T2539;
  wire T2540;
  reg  R2541;
  wire T2542;
  wire T2543;
  wire T2544;
  wire T2545;
  reg [1:0] validVCs_7_2;
  reg  R2546;
  wire T2547;
  wire T2548;
  wire T2549;
  wire T2550;
  reg  R2551;
  wire T2552;
  wire T2553;
  wire T2554;
  wire T2555;
  reg [1:0] validVCs_7_3;
  reg  R2556;
  wire T2557;
  wire T2558;
  wire T2559;
  wire T2560;
  reg  R2561;
  wire T2562;
  wire T2563;
  wire T2564;
  wire T2565;
  reg [1:0] validVCs_7_4;
  reg  R2566;
  wire T2567;
  wire T2568;
  wire T2569;
  wire T2570;
  reg  R2571;
  wire T2572;
  wire T2573;
  wire T2574;
  wire T2575;
  reg [1:0] validVCs_8_0;
  reg  R2576;
  wire T2577;
  wire T2578;
  wire T2579;
  wire T2580;
  reg  R2581;
  wire T2582;
  wire T2583;
  wire T2584;
  wire T2585;
  reg [1:0] validVCs_8_1;
  reg  R2586;
  wire T2587;
  wire T2588;
  wire T2589;
  wire T2590;
  reg  R2591;
  wire T2592;
  wire T2593;
  wire T2594;
  wire T2595;
  reg [1:0] validVCs_8_2;
  reg  R2596;
  wire T2597;
  wire T2598;
  wire T2599;
  wire T2600;
  reg  R2601;
  wire T2602;
  wire T2603;
  wire T2604;
  wire T2605;
  reg [1:0] validVCs_8_3;
  reg  R2606;
  wire T2607;
  wire T2608;
  wire T2609;
  wire T2610;
  reg  R2611;
  wire T2612;
  wire T2613;
  wire T2614;
  wire T2615;
  reg [1:0] validVCs_8_4;
  reg  R2616;
  wire T2617;
  wire T2618;
  wire T2619;
  wire T2620;
  reg  R2621;
  wire T2622;
  wire T2623;
  wire T2624;
  wire T2625;
  reg [1:0] validVCs_9_0;
  reg  R2626;
  wire T2627;
  wire T2628;
  wire T2629;
  wire T2630;
  reg  R2631;
  wire T2632;
  wire T2633;
  wire T2634;
  wire T2635;
  reg [1:0] validVCs_9_1;
  reg  R2636;
  wire T2637;
  wire T2638;
  wire T2639;
  wire T2640;
  reg  R2641;
  wire T2642;
  wire T2643;
  wire T2644;
  wire T2645;
  reg [1:0] validVCs_9_2;
  reg  R2646;
  wire T2647;
  wire T2648;
  wire T2649;
  wire T2650;
  reg  R2651;
  wire T2652;
  wire T2653;
  wire T2654;
  wire T2655;
  reg [1:0] validVCs_9_3;
  reg  R2656;
  wire T2657;
  wire T2658;
  wire T2659;
  wire T2660;
  reg  R2661;
  wire T2662;
  wire T2663;
  wire T2664;
  wire T2665;
  reg [1:0] validVCs_9_4;
  reg  R2666;
  wire T2667;
  wire T2668;
  wire T2669;
  wire T2670;
  reg  R2671;
  wire T2672;
  wire T2673;
  wire T2674;
  reg [2:0] R2675;
  wire[2:0] T3182;
  wire[2:0] T2676;
  wire[2:0] T2677;
  wire[30:0] T2678;
  wire T2679;
  wire T2680;
  wire T2681;
  wire T2682;
  reg [7:0] R2683;
  wire[7:0] T3183;
  wire[7:0] T2684;
  wire T2685;
  wire T2686;
  wire T2687;
  reg  R2688;
  wire T3184;
  reg [2:0] R2689;
  wire[2:0] T3185;
  wire[2:0] T2690;
  wire[2:0] T2691;
  wire[30:0] T2692;
  wire T2693;
  wire T2694;
  wire T2695;
  wire T2696;
  reg [7:0] R2697;
  wire[7:0] T3186;
  wire[7:0] T2698;
  wire T2699;
  wire T2700;
  wire T2701;
  reg  R2702;
  wire T3187;
  reg [2:0] R2703;
  wire[2:0] T3188;
  wire[2:0] T2704;
  wire[2:0] T2705;
  wire[30:0] T2706;
  wire T2707;
  wire T2708;
  wire T2709;
  wire T2710;
  reg [7:0] R2711;
  wire[7:0] T3189;
  wire[7:0] T2712;
  wire T2713;
  wire T2714;
  wire T2715;
  reg  R2716;
  wire T3190;
  reg [2:0] R2717;
  wire[2:0] T3191;
  wire[2:0] T2718;
  wire[2:0] T2719;
  wire[30:0] T2720;
  wire T2721;
  wire T2722;
  wire T2723;
  wire T2724;
  reg [7:0] R2725;
  wire[7:0] T3192;
  wire[7:0] T2726;
  wire T2727;
  wire T2728;
  wire T2729;
  reg  R2730;
  wire T3193;
  reg [2:0] R2731;
  wire[2:0] T3194;
  wire[2:0] T2732;
  wire[2:0] T2733;
  wire[30:0] T2734;
  wire T2735;
  wire T2736;
  wire T2737;
  wire T2738;
  reg [7:0] R2739;
  wire[7:0] T3195;
  wire[7:0] T2740;
  wire T2741;
  wire T2742;
  wire T2743;
  reg  R2744;
  wire T3196;
  reg [2:0] R2745;
  wire[2:0] T3197;
  wire[2:0] T2746;
  wire[2:0] T2747;
  wire[30:0] T2748;
  wire T2749;
  wire T2750;
  wire T2751;
  wire T2752;
  reg [7:0] R2753;
  wire[7:0] T3198;
  wire[7:0] T2754;
  wire T2755;
  wire T2756;
  wire T2757;
  reg  R2758;
  wire T3199;
  reg [2:0] R2759;
  wire[2:0] T3200;
  wire[2:0] T2760;
  wire[2:0] T2761;
  wire[30:0] T2762;
  wire T2763;
  wire T2764;
  wire T2765;
  wire T2766;
  reg [7:0] R2767;
  wire[7:0] T3201;
  wire[7:0] T2768;
  wire T2769;
  wire T2770;
  wire T2771;
  reg  R2772;
  wire T3202;
  reg [2:0] R2773;
  wire[2:0] T3203;
  wire[2:0] T2774;
  wire[2:0] T2775;
  wire[30:0] T2776;
  wire T2777;
  wire T2778;
  wire T2779;
  wire T2780;
  reg [7:0] R2781;
  wire[7:0] T3204;
  wire[7:0] T2782;
  wire T2783;
  wire T2784;
  wire T2785;
  reg  R2786;
  wire T3205;
  reg [2:0] R2787;
  wire[2:0] T3206;
  wire[2:0] T2788;
  wire[2:0] T2789;
  wire[30:0] T2790;
  wire T2791;
  wire T2792;
  wire T2793;
  wire T2794;
  reg [7:0] R2795;
  wire[7:0] T3207;
  wire[7:0] T2796;
  wire T2797;
  wire T2798;
  wire T2799;
  reg  R2800;
  wire T3208;
  reg [2:0] R2801;
  wire[2:0] T3209;
  wire[2:0] T2802;
  wire[2:0] T2803;
  wire[30:0] T2804;
  wire T2805;
  wire T2806;
  wire T2807;
  wire T2808;
  reg [7:0] R2809;
  wire[7:0] T3210;
  wire[7:0] T2810;
  wire T2811;
  wire T2812;
  wire T2813;
  reg  R2814;
  wire T3211;
  wire T2815;
  wire T2816;
  wire T2817;
  wire T2818;
  wire T2819;
  wire T2820;
  wire T2821;
  wire T2822;
  wire T2823;
  wire T2824;
  wire T2825;
  wire T2826;
  wire T2827;
  wire T2828;
  wire T2829;
  wire T2830;
  wire T2831;
  wire T2832;
  wire T2833;
  wire T2834;
  wire T2835;
  wire T2836;
  wire T2837;
  wire T2838;
  wire T2839;
  wire T2840;
  wire T2841;
  wire T2842;
  wire T2843;
  wire T2844;
  wire T2845;
  wire T2846;
  wire T2847;
  wire T2848;
  wire T2849;
  wire T2850;
  wire T2851;
  wire T2852;
  wire T2853;
  wire T2854;
  wire T2855;
  wire T2856;
  wire T2857;
  wire T2858;
  wire T2859;
  wire T2860;
  wire T2861;
  wire T2862;
  wire T2863;
  wire T2864;
  wire T2865;
  wire T2866;
  wire T2867;
  wire T2868;
  wire T2869;
  wire T2870;
  wire T2871;
  wire T2872;
  wire T2873;
  wire T2874;
  wire T2875;
  wire T2876;
  wire T2877;
  wire T2878;
  wire T2879;
  wire T2880;
  wire T2881;
  wire T2882;
  wire T2883;
  wire T2884;
  wire T2885;
  wire T2886;
  wire T2887;
  wire T2888;
  wire T2889;
  wire T2890;
  wire T2891;
  wire T2892;
  wire T2893;
  wire T2894;
  wire T2895;
  wire T2896;
  wire T2897;
  wire T2898;
  wire T2899;
  wire T2900;
  wire T2901;
  wire T2902;
  wire T2903;
  wire T2904;
  wire T2905;
  wire T2906;
  wire T2907;
  wire T2908;
  wire T2909;
  wire T2910;
  wire T2911;
  wire T2912;
  wire T2913;
  wire T2914;
  wire T2915;
  wire T2916;
  wire T2917;
  wire T2918;
  wire T2919;
  wire T2920;
  wire T2921;
  wire T2922;
  wire T2923;
  wire T2924;
  wire T2925;
  wire T2926;
  wire T2927;
  wire T2928;
  wire T2929;
  wire T2930;
  wire T2931;
  wire T2932;
  wire T2933;
  wire T2934;
  wire T2935;
  wire T2936;
  wire T2937;
  wire T2938;
  wire T2939;
  wire T2940;
  wire T2941;
  wire T2942;
  wire T2943;
  wire T2944;
  wire T2945;
  wire T2946;
  wire T2947;
  wire T2948;
  wire T2949;
  wire T2950;
  wire T2951;
  wire T2952;
  wire T2953;
  wire T2954;
  wire T2955;
  wire T2956;
  wire T2957;
  wire T2958;
  wire T2959;
  wire T2960;
  wire T2961;
  wire T2962;
  wire T2963;
  wire T2964;
  wire T2965;
  wire T2966;
  wire T2967;
  wire T2968;
  wire T2969;
  wire T2970;
  wire T2971;
  wire T2972;
  wire T2973;
  wire T2974;
  wire T2975;
  wire T2976;
  wire T2977;
  wire T2978;
  wire T2979;
  wire T2980;
  wire T2981;
  wire T2982;
  wire T2983;
  wire T2984;
  wire T2985;
  wire T2986;
  wire T2987;
  wire T2988;
  wire T2989;
  wire T2990;
  wire T2991;
  wire T2992;
  wire T2993;
  wire T2994;
  wire T2995;
  wire T2996;
  wire T2997;
  wire T2998;
  wire T2999;
  wire T3000;
  wire T3001;
  wire T3002;
  wire T3003;
  wire T3004;
  wire T3005;
  wire T3006;
  wire T3007;
  wire T3008;
  wire T3009;
  wire T3010;
  wire T3011;
  wire T3012;
  wire T3013;
  wire T3014;
  wire T3015;
  wire T3016;
  wire T3017;
  wire T3018;
  wire T3019;
  wire T3020;
  wire T3021;
  wire T3022;
  wire T3023;
  wire T3024;
  wire T3025;
  wire T3026;
  wire T3027;
  wire T3028;
  wire T3029;
  wire T3030;
  wire T3031;
  wire T3032;
  wire T3033;
  wire T3034;
  wire T3035;
  wire T3036;
  wire T3037;
  wire T3038;
  wire T3039;
  wire T3040;
  wire T3041;
  wire T3042;
  wire T3043;
  wire T3044;
  wire T3045;
  wire T3046;
  wire T3047;
  wire T3048;
  wire T3049;
  wire T3050;
  wire T3051;
  wire T3052;
  wire T3053;
  wire T3054;
  wire T3055;
  wire T3056;
  wire T3057;
  wire T3058;
  wire T3059;
  wire T3060;
  wire T3061;
  wire T3062;
  wire T3063;
  wire T3064;
  wire T3065;
  wire T3066;
  wire T3067;
  wire T3068;
  wire T3069;
  wire T3070;
  wire T3071;
  wire T3072;
  wire T3073;
  wire T3074;
  wire T3075;
  wire T3076;
  wire T3077;
  wire T3078;
  wire T3079;
  wire T3080;
  wire T3081;
  wire T3082;
  wire T3083;
  wire T3084;
  wire T3085;
  wire T3086;
  wire T3087;
  wire T3088;
  wire T3089;
  wire T3090;
  wire T3091;
  wire T3092;
  wire T3093;
  wire T3094;
  wire[31:0] T3212;
  wire T3095;
  wire T3096;
  reg  R3097;
  reg [54:0] R3098;
  wire[54:0] T3099;
  wire[54:0] T3213;
  reg  R3100;
  reg [54:0] R3101;
  wire[54:0] T3102;
  wire[54:0] T3214;
  reg  R3103;
  reg [54:0] R3104;
  wire[54:0] T3105;
  wire[54:0] T3215;
  reg  R3106;
  reg [54:0] R3107;
  wire[54:0] T3108;
  wire[54:0] T3216;
  reg  R3109;
  reg [54:0] R3110;
  wire[54:0] T3111;
  wire[54:0] T3217;
  wire[1:0] VCRouterOutputStateManagement_io_currentState;
  wire[1:0] VCRouterOutputStateManagement_1_io_currentState;
  wire[1:0] VCRouterOutputStateManagement_2_io_currentState;
  wire[1:0] VCRouterOutputStateManagement_3_io_currentState;
  wire[1:0] VCRouterOutputStateManagement_4_io_currentState;
  wire CreditGen_io_outCredit_grant;
  wire[54:0] RouterRegFile_io_readData;
  wire RouterRegFile_io_readValid;
  wire[54:0] RouterRegFile_io_readPipelineReg_1;
  wire[54:0] RouterRegFile_io_readPipelineReg_0;
  wire RouterRegFile_io_rvPipelineReg_1;
  wire RouterRegFile_io_rvPipelineReg_0;
  wire[15:0] CMeshDOR_io_outHeadFlit_packetID;
  wire CMeshDOR_io_outHeadFlit_isTail;
  wire CMeshDOR_io_outHeadFlit_vcPort;
  wire[3:0] CMeshDOR_io_outHeadFlit_packetType;
  wire[1:0] CMeshDOR_io_outHeadFlit_destination_2;
  wire[1:0] CMeshDOR_io_outHeadFlit_destination_1;
  wire[1:0] CMeshDOR_io_outHeadFlit_destination_0;
  wire[2:0] CMeshDOR_io_outHeadFlit_priorityLevel;
  wire[2:0] CMeshDOR_io_result;
  wire[1:0] CMeshDOR_io_vcsAvailable_4;
  wire[1:0] CMeshDOR_io_vcsAvailable_3;
  wire[1:0] CMeshDOR_io_vcsAvailable_2;
  wire[1:0] CMeshDOR_io_vcsAvailable_1;
  wire[1:0] CMeshDOR_io_vcsAvailable_0;
  wire[2:0] VCRouterStateManagement_io_currentState;
  wire CreditGen_1_io_outCredit_grant;
  wire[54:0] RouterRegFile_1_io_readData;
  wire RouterRegFile_1_io_readValid;
  wire[54:0] RouterRegFile_1_io_readPipelineReg_1;
  wire[54:0] RouterRegFile_1_io_readPipelineReg_0;
  wire RouterRegFile_1_io_rvPipelineReg_1;
  wire RouterRegFile_1_io_rvPipelineReg_0;
  wire[15:0] CMeshDOR_1_io_outHeadFlit_packetID;
  wire CMeshDOR_1_io_outHeadFlit_isTail;
  wire CMeshDOR_1_io_outHeadFlit_vcPort;
  wire[3:0] CMeshDOR_1_io_outHeadFlit_packetType;
  wire[1:0] CMeshDOR_1_io_outHeadFlit_destination_2;
  wire[1:0] CMeshDOR_1_io_outHeadFlit_destination_1;
  wire[1:0] CMeshDOR_1_io_outHeadFlit_destination_0;
  wire[2:0] CMeshDOR_1_io_outHeadFlit_priorityLevel;
  wire[2:0] CMeshDOR_1_io_result;
  wire[1:0] CMeshDOR_1_io_vcsAvailable_4;
  wire[1:0] CMeshDOR_1_io_vcsAvailable_3;
  wire[1:0] CMeshDOR_1_io_vcsAvailable_2;
  wire[1:0] CMeshDOR_1_io_vcsAvailable_1;
  wire[1:0] CMeshDOR_1_io_vcsAvailable_0;
  wire[2:0] VCRouterStateManagement_1_io_currentState;
  wire CreditGen_2_io_outCredit_grant;
  wire[54:0] RouterRegFile_2_io_readData;
  wire RouterRegFile_2_io_readValid;
  wire[54:0] RouterRegFile_2_io_readPipelineReg_1;
  wire[54:0] RouterRegFile_2_io_readPipelineReg_0;
  wire RouterRegFile_2_io_rvPipelineReg_1;
  wire RouterRegFile_2_io_rvPipelineReg_0;
  wire[15:0] CMeshDOR_2_io_outHeadFlit_packetID;
  wire CMeshDOR_2_io_outHeadFlit_isTail;
  wire CMeshDOR_2_io_outHeadFlit_vcPort;
  wire[3:0] CMeshDOR_2_io_outHeadFlit_packetType;
  wire[1:0] CMeshDOR_2_io_outHeadFlit_destination_2;
  wire[1:0] CMeshDOR_2_io_outHeadFlit_destination_1;
  wire[1:0] CMeshDOR_2_io_outHeadFlit_destination_0;
  wire[2:0] CMeshDOR_2_io_outHeadFlit_priorityLevel;
  wire[2:0] CMeshDOR_2_io_result;
  wire[1:0] CMeshDOR_2_io_vcsAvailable_4;
  wire[1:0] CMeshDOR_2_io_vcsAvailable_3;
  wire[1:0] CMeshDOR_2_io_vcsAvailable_2;
  wire[1:0] CMeshDOR_2_io_vcsAvailable_1;
  wire[1:0] CMeshDOR_2_io_vcsAvailable_0;
  wire[2:0] VCRouterStateManagement_2_io_currentState;
  wire CreditGen_3_io_outCredit_grant;
  wire[54:0] RouterRegFile_3_io_readData;
  wire RouterRegFile_3_io_readValid;
  wire[54:0] RouterRegFile_3_io_readPipelineReg_1;
  wire[54:0] RouterRegFile_3_io_readPipelineReg_0;
  wire RouterRegFile_3_io_rvPipelineReg_1;
  wire RouterRegFile_3_io_rvPipelineReg_0;
  wire[15:0] CMeshDOR_3_io_outHeadFlit_packetID;
  wire CMeshDOR_3_io_outHeadFlit_isTail;
  wire CMeshDOR_3_io_outHeadFlit_vcPort;
  wire[3:0] CMeshDOR_3_io_outHeadFlit_packetType;
  wire[1:0] CMeshDOR_3_io_outHeadFlit_destination_2;
  wire[1:0] CMeshDOR_3_io_outHeadFlit_destination_1;
  wire[1:0] CMeshDOR_3_io_outHeadFlit_destination_0;
  wire[2:0] CMeshDOR_3_io_outHeadFlit_priorityLevel;
  wire[2:0] CMeshDOR_3_io_result;
  wire[1:0] CMeshDOR_3_io_vcsAvailable_4;
  wire[1:0] CMeshDOR_3_io_vcsAvailable_3;
  wire[1:0] CMeshDOR_3_io_vcsAvailable_2;
  wire[1:0] CMeshDOR_3_io_vcsAvailable_1;
  wire[1:0] CMeshDOR_3_io_vcsAvailable_0;
  wire[2:0] VCRouterStateManagement_3_io_currentState;
  wire CreditGen_4_io_outCredit_grant;
  wire[54:0] RouterRegFile_4_io_readData;
  wire RouterRegFile_4_io_readValid;
  wire[54:0] RouterRegFile_4_io_readPipelineReg_1;
  wire[54:0] RouterRegFile_4_io_readPipelineReg_0;
  wire RouterRegFile_4_io_rvPipelineReg_1;
  wire RouterRegFile_4_io_rvPipelineReg_0;
  wire[15:0] CMeshDOR_4_io_outHeadFlit_packetID;
  wire CMeshDOR_4_io_outHeadFlit_isTail;
  wire CMeshDOR_4_io_outHeadFlit_vcPort;
  wire[3:0] CMeshDOR_4_io_outHeadFlit_packetType;
  wire[1:0] CMeshDOR_4_io_outHeadFlit_destination_2;
  wire[1:0] CMeshDOR_4_io_outHeadFlit_destination_1;
  wire[1:0] CMeshDOR_4_io_outHeadFlit_destination_0;
  wire[2:0] CMeshDOR_4_io_outHeadFlit_priorityLevel;
  wire[2:0] CMeshDOR_4_io_result;
  wire[1:0] CMeshDOR_4_io_vcsAvailable_4;
  wire[1:0] CMeshDOR_4_io_vcsAvailable_3;
  wire[1:0] CMeshDOR_4_io_vcsAvailable_2;
  wire[1:0] CMeshDOR_4_io_vcsAvailable_1;
  wire[1:0] CMeshDOR_4_io_vcsAvailable_0;
  wire[2:0] VCRouterStateManagement_4_io_currentState;
  wire CreditGen_5_io_outCredit_grant;
  wire[54:0] RouterRegFile_5_io_readData;
  wire RouterRegFile_5_io_readValid;
  wire[54:0] RouterRegFile_5_io_readPipelineReg_1;
  wire[54:0] RouterRegFile_5_io_readPipelineReg_0;
  wire RouterRegFile_5_io_rvPipelineReg_1;
  wire RouterRegFile_5_io_rvPipelineReg_0;
  wire[15:0] CMeshDOR_5_io_outHeadFlit_packetID;
  wire CMeshDOR_5_io_outHeadFlit_isTail;
  wire CMeshDOR_5_io_outHeadFlit_vcPort;
  wire[3:0] CMeshDOR_5_io_outHeadFlit_packetType;
  wire[1:0] CMeshDOR_5_io_outHeadFlit_destination_2;
  wire[1:0] CMeshDOR_5_io_outHeadFlit_destination_1;
  wire[1:0] CMeshDOR_5_io_outHeadFlit_destination_0;
  wire[2:0] CMeshDOR_5_io_outHeadFlit_priorityLevel;
  wire[2:0] CMeshDOR_5_io_result;
  wire[1:0] CMeshDOR_5_io_vcsAvailable_4;
  wire[1:0] CMeshDOR_5_io_vcsAvailable_3;
  wire[1:0] CMeshDOR_5_io_vcsAvailable_2;
  wire[1:0] CMeshDOR_5_io_vcsAvailable_1;
  wire[1:0] CMeshDOR_5_io_vcsAvailable_0;
  wire[2:0] VCRouterStateManagement_5_io_currentState;
  wire CreditGen_6_io_outCredit_grant;
  wire[54:0] RouterRegFile_6_io_readData;
  wire RouterRegFile_6_io_readValid;
  wire[54:0] RouterRegFile_6_io_readPipelineReg_1;
  wire[54:0] RouterRegFile_6_io_readPipelineReg_0;
  wire RouterRegFile_6_io_rvPipelineReg_1;
  wire RouterRegFile_6_io_rvPipelineReg_0;
  wire[15:0] CMeshDOR_6_io_outHeadFlit_packetID;
  wire CMeshDOR_6_io_outHeadFlit_isTail;
  wire CMeshDOR_6_io_outHeadFlit_vcPort;
  wire[3:0] CMeshDOR_6_io_outHeadFlit_packetType;
  wire[1:0] CMeshDOR_6_io_outHeadFlit_destination_2;
  wire[1:0] CMeshDOR_6_io_outHeadFlit_destination_1;
  wire[1:0] CMeshDOR_6_io_outHeadFlit_destination_0;
  wire[2:0] CMeshDOR_6_io_outHeadFlit_priorityLevel;
  wire[2:0] CMeshDOR_6_io_result;
  wire[1:0] CMeshDOR_6_io_vcsAvailable_4;
  wire[1:0] CMeshDOR_6_io_vcsAvailable_3;
  wire[1:0] CMeshDOR_6_io_vcsAvailable_2;
  wire[1:0] CMeshDOR_6_io_vcsAvailable_1;
  wire[1:0] CMeshDOR_6_io_vcsAvailable_0;
  wire[2:0] VCRouterStateManagement_6_io_currentState;
  wire CreditGen_7_io_outCredit_grant;
  wire[54:0] RouterRegFile_7_io_readData;
  wire RouterRegFile_7_io_readValid;
  wire[54:0] RouterRegFile_7_io_readPipelineReg_1;
  wire[54:0] RouterRegFile_7_io_readPipelineReg_0;
  wire RouterRegFile_7_io_rvPipelineReg_1;
  wire RouterRegFile_7_io_rvPipelineReg_0;
  wire[15:0] CMeshDOR_7_io_outHeadFlit_packetID;
  wire CMeshDOR_7_io_outHeadFlit_isTail;
  wire CMeshDOR_7_io_outHeadFlit_vcPort;
  wire[3:0] CMeshDOR_7_io_outHeadFlit_packetType;
  wire[1:0] CMeshDOR_7_io_outHeadFlit_destination_2;
  wire[1:0] CMeshDOR_7_io_outHeadFlit_destination_1;
  wire[1:0] CMeshDOR_7_io_outHeadFlit_destination_0;
  wire[2:0] CMeshDOR_7_io_outHeadFlit_priorityLevel;
  wire[2:0] CMeshDOR_7_io_result;
  wire[1:0] CMeshDOR_7_io_vcsAvailable_4;
  wire[1:0] CMeshDOR_7_io_vcsAvailable_3;
  wire[1:0] CMeshDOR_7_io_vcsAvailable_2;
  wire[1:0] CMeshDOR_7_io_vcsAvailable_1;
  wire[1:0] CMeshDOR_7_io_vcsAvailable_0;
  wire[2:0] VCRouterStateManagement_7_io_currentState;
  wire CreditGen_8_io_outCredit_grant;
  wire[54:0] RouterRegFile_8_io_readData;
  wire RouterRegFile_8_io_readValid;
  wire[54:0] RouterRegFile_8_io_readPipelineReg_1;
  wire[54:0] RouterRegFile_8_io_readPipelineReg_0;
  wire RouterRegFile_8_io_rvPipelineReg_1;
  wire RouterRegFile_8_io_rvPipelineReg_0;
  wire[15:0] CMeshDOR_8_io_outHeadFlit_packetID;
  wire CMeshDOR_8_io_outHeadFlit_isTail;
  wire CMeshDOR_8_io_outHeadFlit_vcPort;
  wire[3:0] CMeshDOR_8_io_outHeadFlit_packetType;
  wire[1:0] CMeshDOR_8_io_outHeadFlit_destination_2;
  wire[1:0] CMeshDOR_8_io_outHeadFlit_destination_1;
  wire[1:0] CMeshDOR_8_io_outHeadFlit_destination_0;
  wire[2:0] CMeshDOR_8_io_outHeadFlit_priorityLevel;
  wire[2:0] CMeshDOR_8_io_result;
  wire[1:0] CMeshDOR_8_io_vcsAvailable_4;
  wire[1:0] CMeshDOR_8_io_vcsAvailable_3;
  wire[1:0] CMeshDOR_8_io_vcsAvailable_2;
  wire[1:0] CMeshDOR_8_io_vcsAvailable_1;
  wire[1:0] CMeshDOR_8_io_vcsAvailable_0;
  wire[2:0] VCRouterStateManagement_8_io_currentState;
  wire CreditGen_9_io_outCredit_grant;
  wire[54:0] RouterRegFile_9_io_readData;
  wire RouterRegFile_9_io_readValid;
  wire[54:0] RouterRegFile_9_io_readPipelineReg_1;
  wire[54:0] RouterRegFile_9_io_readPipelineReg_0;
  wire RouterRegFile_9_io_rvPipelineReg_1;
  wire RouterRegFile_9_io_rvPipelineReg_0;
  wire[15:0] CMeshDOR_9_io_outHeadFlit_packetID;
  wire CMeshDOR_9_io_outHeadFlit_isTail;
  wire CMeshDOR_9_io_outHeadFlit_vcPort;
  wire[3:0] CMeshDOR_9_io_outHeadFlit_packetType;
  wire[1:0] CMeshDOR_9_io_outHeadFlit_destination_2;
  wire[1:0] CMeshDOR_9_io_outHeadFlit_destination_1;
  wire[1:0] CMeshDOR_9_io_outHeadFlit_destination_0;
  wire[2:0] CMeshDOR_9_io_outHeadFlit_priorityLevel;
  wire[2:0] CMeshDOR_9_io_result;
  wire[1:0] CMeshDOR_9_io_vcsAvailable_4;
  wire[1:0] CMeshDOR_9_io_vcsAvailable_3;
  wire[1:0] CMeshDOR_9_io_vcsAvailable_2;
  wire[1:0] CMeshDOR_9_io_vcsAvailable_1;
  wire[1:0] CMeshDOR_9_io_vcsAvailable_0;
  wire[2:0] VCRouterStateManagement_9_io_currentState;
  wire CreditCon_io_outCredit;
  wire CreditCon_1_io_outCredit;
  wire CreditCon_2_io_outCredit;
  wire CreditCon_3_io_outCredit;
  wire CreditCon_4_io_outCredit;
  wire CreditCon_5_io_outCredit;
  wire CreditCon_6_io_outCredit;
  wire CreditCon_7_io_outCredit;
  wire CreditCon_8_io_outCredit;
  wire CreditCon_9_io_outCredit;
  wire[54:0] switch_io_outPorts_4_x;
  wire[54:0] switch_io_outPorts_3_x;
  wire[54:0] switch_io_outPorts_2_x;
  wire[54:0] switch_io_outPorts_1_x;
  wire[54:0] switch_io_outPorts_0_x;
  wire swAllocator_io_requests_4_9_grant;
  wire swAllocator_io_requests_4_8_grant;
  wire swAllocator_io_requests_4_7_grant;
  wire swAllocator_io_requests_4_6_grant;
  wire swAllocator_io_requests_4_5_grant;
  wire swAllocator_io_requests_4_4_grant;
  wire swAllocator_io_requests_4_3_grant;
  wire swAllocator_io_requests_4_2_grant;
  wire swAllocator_io_requests_4_1_grant;
  wire swAllocator_io_requests_4_0_grant;
  wire swAllocator_io_requests_3_9_grant;
  wire swAllocator_io_requests_3_8_grant;
  wire swAllocator_io_requests_3_7_grant;
  wire swAllocator_io_requests_3_6_grant;
  wire swAllocator_io_requests_3_5_grant;
  wire swAllocator_io_requests_3_4_grant;
  wire swAllocator_io_requests_3_3_grant;
  wire swAllocator_io_requests_3_2_grant;
  wire swAllocator_io_requests_3_1_grant;
  wire swAllocator_io_requests_3_0_grant;
  wire swAllocator_io_requests_2_9_grant;
  wire swAllocator_io_requests_2_8_grant;
  wire swAllocator_io_requests_2_7_grant;
  wire swAllocator_io_requests_2_6_grant;
  wire swAllocator_io_requests_2_5_grant;
  wire swAllocator_io_requests_2_4_grant;
  wire swAllocator_io_requests_2_3_grant;
  wire swAllocator_io_requests_2_2_grant;
  wire swAllocator_io_requests_2_1_grant;
  wire swAllocator_io_requests_2_0_grant;
  wire swAllocator_io_requests_1_9_grant;
  wire swAllocator_io_requests_1_8_grant;
  wire swAllocator_io_requests_1_7_grant;
  wire swAllocator_io_requests_1_6_grant;
  wire swAllocator_io_requests_1_5_grant;
  wire swAllocator_io_requests_1_4_grant;
  wire swAllocator_io_requests_1_3_grant;
  wire swAllocator_io_requests_1_2_grant;
  wire swAllocator_io_requests_1_1_grant;
  wire swAllocator_io_requests_1_0_grant;
  wire swAllocator_io_requests_0_9_grant;
  wire swAllocator_io_requests_0_8_grant;
  wire swAllocator_io_requests_0_7_grant;
  wire swAllocator_io_requests_0_6_grant;
  wire swAllocator_io_requests_0_5_grant;
  wire swAllocator_io_requests_0_4_grant;
  wire swAllocator_io_requests_0_3_grant;
  wire swAllocator_io_requests_0_2_grant;
  wire swAllocator_io_requests_0_1_grant;
  wire swAllocator_io_requests_0_0_grant;
  wire[3:0] swAllocator_io_chosens_4;
  wire[3:0] swAllocator_io_chosens_3;
  wire[3:0] swAllocator_io_chosens_2;
  wire[3:0] swAllocator_io_chosens_1;
  wire[3:0] swAllocator_io_chosens_0;
  wire vcAllocator_io_resources_9_valid;
  wire vcAllocator_io_resources_8_valid;
  wire vcAllocator_io_resources_7_valid;
  wire vcAllocator_io_resources_6_valid;
  wire vcAllocator_io_resources_5_valid;
  wire vcAllocator_io_resources_4_valid;
  wire vcAllocator_io_resources_3_valid;
  wire vcAllocator_io_resources_2_valid;
  wire vcAllocator_io_resources_1_valid;
  wire vcAllocator_io_resources_0_valid;
  wire[3:0] vcAllocator_io_chosens_9;
  wire[3:0] vcAllocator_io_chosens_8;
  wire[3:0] vcAllocator_io_chosens_7;
  wire[3:0] vcAllocator_io_chosens_6;
  wire[3:0] vcAllocator_io_chosens_5;
  wire[3:0] vcAllocator_io_chosens_4;
  wire[3:0] vcAllocator_io_chosens_3;
  wire[3:0] vcAllocator_io_chosens_2;
  wire[3:0] vcAllocator_io_chosens_1;
  wire[3:0] vcAllocator_io_chosens_0;
  wire RouterBuffer_io_enq_ready;
  wire RouterBuffer_io_deq_valid;
  wire[54:0] RouterBuffer_io_deq_bits_x;
  wire[54:0] ReplaceVCPort_io_newFlit_x;
  wire RouterBuffer_1_io_enq_ready;
  wire RouterBuffer_1_io_deq_valid;
  wire[54:0] RouterBuffer_1_io_deq_bits_x;
  wire[54:0] ReplaceVCPort_1_io_newFlit_x;
  wire RouterBuffer_2_io_enq_ready;
  wire RouterBuffer_2_io_deq_valid;
  wire[54:0] RouterBuffer_2_io_deq_bits_x;
  wire[54:0] ReplaceVCPort_2_io_newFlit_x;
  wire RouterBuffer_3_io_enq_ready;
  wire RouterBuffer_3_io_deq_valid;
  wire[54:0] RouterBuffer_3_io_deq_bits_x;
  wire[54:0] ReplaceVCPort_3_io_newFlit_x;
  wire RouterBuffer_4_io_enq_ready;
  wire RouterBuffer_4_io_deq_valid;
  wire[54:0] RouterBuffer_4_io_deq_bits_x;
  wire[54:0] ReplaceVCPort_4_io_newFlit_x;
  wire RouterBuffer_5_io_enq_ready;
  wire RouterBuffer_5_io_deq_valid;
  wire[54:0] RouterBuffer_5_io_deq_bits_x;
  wire[54:0] ReplaceVCPort_5_io_newFlit_x;
  wire RouterBuffer_6_io_enq_ready;
  wire RouterBuffer_6_io_deq_valid;
  wire[54:0] RouterBuffer_6_io_deq_bits_x;
  wire[54:0] ReplaceVCPort_6_io_newFlit_x;
  wire RouterBuffer_7_io_enq_ready;
  wire RouterBuffer_7_io_deq_valid;
  wire[54:0] RouterBuffer_7_io_deq_bits_x;
  wire[54:0] ReplaceVCPort_7_io_newFlit_x;
  wire RouterBuffer_8_io_enq_ready;
  wire RouterBuffer_8_io_deq_valid;
  wire[54:0] RouterBuffer_8_io_deq_bits_x;
  wire[54:0] ReplaceVCPort_8_io_newFlit_x;
  wire RouterBuffer_9_io_enq_ready;
  wire RouterBuffer_9_io_deq_valid;
  wire[54:0] RouterBuffer_9_io_deq_bits_x;
  wire[54:0] ReplaceVCPort_9_io_newFlit_x;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    T0 = 1'b0;
    T17 = 1'b0;
    T22 = 1'b0;
    T39 = 1'b0;
    T44 = 1'b0;
    T61 = 1'b0;
    T66 = 1'b0;
    T83 = 1'b0;
    T88 = 1'b0;
    T105 = 1'b0;
    T110 = 1'b0;
    T127 = 1'b0;
    T132 = 1'b0;
    T149 = 1'b0;
    T154 = 1'b0;
    T171 = 1'b0;
    T176 = 1'b0;
    T193 = 1'b0;
    T198 = 1'b0;
    T215 = 1'b0;
    R282 = {2{1'b0}};
    R295 = {1{1'b0}};
    R349 = {1{1'b0}};
    R426 = {2{1'b0}};
    R439 = {1{1'b0}};
    R493 = {1{1'b0}};
    R570 = {2{1'b0}};
    R583 = {1{1'b0}};
    R637 = {1{1'b0}};
    R714 = {2{1'b0}};
    R727 = {1{1'b0}};
    R781 = {1{1'b0}};
    R858 = {2{1'b0}};
    R871 = {1{1'b0}};
    R925 = {1{1'b0}};
    R1002 = {2{1'b0}};
    R1015 = {1{1'b0}};
    R1069 = {1{1'b0}};
    R1146 = {2{1'b0}};
    R1159 = {1{1'b0}};
    R1213 = {1{1'b0}};
    R1290 = {2{1'b0}};
    R1303 = {1{1'b0}};
    R1357 = {1{1'b0}};
    R1434 = {2{1'b0}};
    R1447 = {1{1'b0}};
    R1501 = {1{1'b0}};
    R1578 = {2{1'b0}};
    R1591 = {1{1'b0}};
    R1645 = {1{1'b0}};
    validVCs_0_0 = {1{1'b0}};
    R2176 = {1{1'b0}};
    R2181 = {1{1'b0}};
    validVCs_0_1 = {1{1'b0}};
    R2186 = {1{1'b0}};
    R2191 = {1{1'b0}};
    validVCs_0_2 = {1{1'b0}};
    R2196 = {1{1'b0}};
    R2201 = {1{1'b0}};
    validVCs_0_3 = {1{1'b0}};
    R2206 = {1{1'b0}};
    R2211 = {1{1'b0}};
    validVCs_0_4 = {1{1'b0}};
    R2216 = {1{1'b0}};
    R2221 = {1{1'b0}};
    validVCs_1_0 = {1{1'b0}};
    R2226 = {1{1'b0}};
    R2231 = {1{1'b0}};
    validVCs_1_1 = {1{1'b0}};
    R2236 = {1{1'b0}};
    R2241 = {1{1'b0}};
    validVCs_1_2 = {1{1'b0}};
    R2246 = {1{1'b0}};
    R2251 = {1{1'b0}};
    validVCs_1_3 = {1{1'b0}};
    R2256 = {1{1'b0}};
    R2261 = {1{1'b0}};
    validVCs_1_4 = {1{1'b0}};
    R2266 = {1{1'b0}};
    R2271 = {1{1'b0}};
    validVCs_2_0 = {1{1'b0}};
    R2276 = {1{1'b0}};
    R2281 = {1{1'b0}};
    validVCs_2_1 = {1{1'b0}};
    R2286 = {1{1'b0}};
    R2291 = {1{1'b0}};
    validVCs_2_2 = {1{1'b0}};
    R2296 = {1{1'b0}};
    R2301 = {1{1'b0}};
    validVCs_2_3 = {1{1'b0}};
    R2306 = {1{1'b0}};
    R2311 = {1{1'b0}};
    validVCs_2_4 = {1{1'b0}};
    R2316 = {1{1'b0}};
    R2321 = {1{1'b0}};
    validVCs_3_0 = {1{1'b0}};
    R2326 = {1{1'b0}};
    R2331 = {1{1'b0}};
    validVCs_3_1 = {1{1'b0}};
    R2336 = {1{1'b0}};
    R2341 = {1{1'b0}};
    validVCs_3_2 = {1{1'b0}};
    R2346 = {1{1'b0}};
    R2351 = {1{1'b0}};
    validVCs_3_3 = {1{1'b0}};
    R2356 = {1{1'b0}};
    R2361 = {1{1'b0}};
    validVCs_3_4 = {1{1'b0}};
    R2366 = {1{1'b0}};
    R2371 = {1{1'b0}};
    validVCs_4_0 = {1{1'b0}};
    R2376 = {1{1'b0}};
    R2381 = {1{1'b0}};
    validVCs_4_1 = {1{1'b0}};
    R2386 = {1{1'b0}};
    R2391 = {1{1'b0}};
    validVCs_4_2 = {1{1'b0}};
    R2396 = {1{1'b0}};
    R2401 = {1{1'b0}};
    validVCs_4_3 = {1{1'b0}};
    R2406 = {1{1'b0}};
    R2411 = {1{1'b0}};
    validVCs_4_4 = {1{1'b0}};
    R2416 = {1{1'b0}};
    R2421 = {1{1'b0}};
    validVCs_5_0 = {1{1'b0}};
    R2426 = {1{1'b0}};
    R2431 = {1{1'b0}};
    validVCs_5_1 = {1{1'b0}};
    R2436 = {1{1'b0}};
    R2441 = {1{1'b0}};
    validVCs_5_2 = {1{1'b0}};
    R2446 = {1{1'b0}};
    R2451 = {1{1'b0}};
    validVCs_5_3 = {1{1'b0}};
    R2456 = {1{1'b0}};
    R2461 = {1{1'b0}};
    validVCs_5_4 = {1{1'b0}};
    R2466 = {1{1'b0}};
    R2471 = {1{1'b0}};
    validVCs_6_0 = {1{1'b0}};
    R2476 = {1{1'b0}};
    R2481 = {1{1'b0}};
    validVCs_6_1 = {1{1'b0}};
    R2486 = {1{1'b0}};
    R2491 = {1{1'b0}};
    validVCs_6_2 = {1{1'b0}};
    R2496 = {1{1'b0}};
    R2501 = {1{1'b0}};
    validVCs_6_3 = {1{1'b0}};
    R2506 = {1{1'b0}};
    R2511 = {1{1'b0}};
    validVCs_6_4 = {1{1'b0}};
    R2516 = {1{1'b0}};
    R2521 = {1{1'b0}};
    validVCs_7_0 = {1{1'b0}};
    R2526 = {1{1'b0}};
    R2531 = {1{1'b0}};
    validVCs_7_1 = {1{1'b0}};
    R2536 = {1{1'b0}};
    R2541 = {1{1'b0}};
    validVCs_7_2 = {1{1'b0}};
    R2546 = {1{1'b0}};
    R2551 = {1{1'b0}};
    validVCs_7_3 = {1{1'b0}};
    R2556 = {1{1'b0}};
    R2561 = {1{1'b0}};
    validVCs_7_4 = {1{1'b0}};
    R2566 = {1{1'b0}};
    R2571 = {1{1'b0}};
    validVCs_8_0 = {1{1'b0}};
    R2576 = {1{1'b0}};
    R2581 = {1{1'b0}};
    validVCs_8_1 = {1{1'b0}};
    R2586 = {1{1'b0}};
    R2591 = {1{1'b0}};
    validVCs_8_2 = {1{1'b0}};
    R2596 = {1{1'b0}};
    R2601 = {1{1'b0}};
    validVCs_8_3 = {1{1'b0}};
    R2606 = {1{1'b0}};
    R2611 = {1{1'b0}};
    validVCs_8_4 = {1{1'b0}};
    R2616 = {1{1'b0}};
    R2621 = {1{1'b0}};
    validVCs_9_0 = {1{1'b0}};
    R2626 = {1{1'b0}};
    R2631 = {1{1'b0}};
    validVCs_9_1 = {1{1'b0}};
    R2636 = {1{1'b0}};
    R2641 = {1{1'b0}};
    validVCs_9_2 = {1{1'b0}};
    R2646 = {1{1'b0}};
    R2651 = {1{1'b0}};
    validVCs_9_3 = {1{1'b0}};
    R2656 = {1{1'b0}};
    R2661 = {1{1'b0}};
    validVCs_9_4 = {1{1'b0}};
    R2666 = {1{1'b0}};
    R2671 = {1{1'b0}};
    R2675 = {1{1'b0}};
    R2683 = {1{1'b0}};
    R2688 = {1{1'b0}};
    R2689 = {1{1'b0}};
    R2697 = {1{1'b0}};
    R2702 = {1{1'b0}};
    R2703 = {1{1'b0}};
    R2711 = {1{1'b0}};
    R2716 = {1{1'b0}};
    R2717 = {1{1'b0}};
    R2725 = {1{1'b0}};
    R2730 = {1{1'b0}};
    R2731 = {1{1'b0}};
    R2739 = {1{1'b0}};
    R2744 = {1{1'b0}};
    R2745 = {1{1'b0}};
    R2753 = {1{1'b0}};
    R2758 = {1{1'b0}};
    R2759 = {1{1'b0}};
    R2767 = {1{1'b0}};
    R2772 = {1{1'b0}};
    R2773 = {1{1'b0}};
    R2781 = {1{1'b0}};
    R2786 = {1{1'b0}};
    R2787 = {1{1'b0}};
    R2795 = {1{1'b0}};
    R2800 = {1{1'b0}};
    R2801 = {1{1'b0}};
    R2809 = {1{1'b0}};
    R2814 = {1{1'b0}};
    R3097 = {1{1'b0}};
    R3098 = {2{1'b0}};
    R3100 = {1{1'b0}};
    R3101 = {2{1'b0}};
    R3103 = {1{1'b0}};
    R3104 = {2{1'b0}};
    R3106 = {1{1'b0}};
    R3107 = {2{1'b0}};
    R3109 = {1{1'b0}};
    R3110 = {2{1'b0}};
  end
// synthesis translate_on
`endif

`ifndef SYNTHESIS
// synthesis translate_off
//  assign io_counters_0_counterIndex = {1{1'b0}};
//  assign io_counters_1_counterIndex = {1{1'b0}};
//  assign io_counters_1_counterVal = {1{1'b0}};
// synthesis translate_on
`endif
  assign T1 = T2 | reset;
  assign T2 = T13 | T3;
  assign T3 = ~ T4;
  assign T4 = T5 == 1'h1;
  assign T5 = T6;
  assign T6 = T11 ? T9 : T7;
  assign T7 = T8[6'h24:6'h24];
  assign T8 = io_inChannels_4_flit_x[6'h36:1'h1];
  assign T9 = T10[4'hd:4'hd];
  assign T10 = io_inChannels_4_flit_x[5'h1f:1'h1];
  assign T11 = T12 == 1'h1;
  assign T12 = io_inChannels_4_flit_x[1'h0:1'h0];
  assign T13 = T15 | T14;
  assign T14 = ~ io_inChannels_4_flitValid;
  assign T15 = T16 & T4;
  assign T16 = RouterBuffer_9_io_enq_ready & io_inChannels_4_flitValid;
  assign T18 = T19 | reset;
  assign T19 = T21 | T20;
  assign T20 = T379 & T4;
  assign T21 = ~ T379;
  assign T23 = T24 | reset;
  assign T24 = T35 | T25;
  assign T25 = ~ T26;
  assign T26 = T27 == 1'h0;
  assign T27 = T28;
  assign T28 = T33 ? T31 : T29;
  assign T29 = T30[6'h24:6'h24];
  assign T30 = io_inChannels_4_flit_x[6'h36:1'h1];
  assign T31 = T32[4'hd:4'hd];
  assign T32 = io_inChannels_4_flit_x[5'h1f:1'h1];
  assign T33 = T34 == 1'h1;
  assign T34 = io_inChannels_4_flit_x[1'h0:1'h0];
  assign T35 = T37 | T36;
  assign T36 = ~ io_inChannels_4_flitValid;
  assign T37 = T38 & T26;
  assign T38 = RouterBuffer_8_io_enq_ready & io_inChannels_4_flitValid;
  assign T40 = T41 | reset;
  assign T41 = T43 | T42;
  assign T42 = T523 & T26;
  assign T43 = ~ T523;
  assign T45 = T46 | reset;
  assign T46 = T57 | T47;
  assign T47 = ~ T48;
  assign T48 = T49 == 1'h1;
  assign T49 = T50;
  assign T50 = T55 ? T53 : T51;
  assign T51 = T52[6'h24:6'h24];
  assign T52 = io_inChannels_3_flit_x[6'h36:1'h1];
  assign T53 = T54[4'hd:4'hd];
  assign T54 = io_inChannels_3_flit_x[5'h1f:1'h1];
  assign T55 = T56 == 1'h1;
  assign T56 = io_inChannels_3_flit_x[1'h0:1'h0];
  assign T57 = T59 | T58;
  assign T58 = ~ io_inChannels_3_flitValid;
  assign T59 = T60 & T48;
  assign T60 = RouterBuffer_7_io_enq_ready & io_inChannels_3_flitValid;
  assign T62 = T63 | reset;
  assign T63 = T65 | T64;
  assign T64 = T667 & T48;
  assign T65 = ~ T667;
  assign T67 = T68 | reset;
  assign T68 = T79 | T69;
  assign T69 = ~ T70;
  assign T70 = T71 == 1'h0;
  assign T71 = T72;
  assign T72 = T77 ? T75 : T73;
  assign T73 = T74[6'h24:6'h24];
  assign T74 = io_inChannels_3_flit_x[6'h36:1'h1];
  assign T75 = T76[4'hd:4'hd];
  assign T76 = io_inChannels_3_flit_x[5'h1f:1'h1];
  assign T77 = T78 == 1'h1;
  assign T78 = io_inChannels_3_flit_x[1'h0:1'h0];
  assign T79 = T81 | T80;
  assign T80 = ~ io_inChannels_3_flitValid;
  assign T81 = T82 & T70;
  assign T82 = RouterBuffer_6_io_enq_ready & io_inChannels_3_flitValid;
  assign T84 = T85 | reset;
  assign T85 = T87 | T86;
  assign T86 = T811 & T70;
  assign T87 = ~ T811;
  assign T89 = T90 | reset;
  assign T90 = T101 | T91;
  assign T91 = ~ T92;
  assign T92 = T93 == 1'h1;
  assign T93 = T94;
  assign T94 = T99 ? T97 : T95;
  assign T95 = T96[6'h24:6'h24];
  assign T96 = io_inChannels_2_flit_x[6'h36:1'h1];
  assign T97 = T98[4'hd:4'hd];
  assign T98 = io_inChannels_2_flit_x[5'h1f:1'h1];
  assign T99 = T100 == 1'h1;
  assign T100 = io_inChannels_2_flit_x[1'h0:1'h0];
  assign T101 = T103 | T102;
  assign T102 = ~ io_inChannels_2_flitValid;
  assign T103 = T104 & T92;
  assign T104 = RouterBuffer_5_io_enq_ready & io_inChannels_2_flitValid;
  assign T106 = T107 | reset;
  assign T107 = T109 | T108;
  assign T108 = T955 & T92;
  assign T109 = ~ T955;
  assign T111 = T112 | reset;
  assign T112 = T123 | T113;
  assign T113 = ~ T114;
  assign T114 = T115 == 1'h0;
  assign T115 = T116;
  assign T116 = T121 ? T119 : T117;
  assign T117 = T118[6'h24:6'h24];
  assign T118 = io_inChannels_2_flit_x[6'h36:1'h1];
  assign T119 = T120[4'hd:4'hd];
  assign T120 = io_inChannels_2_flit_x[5'h1f:1'h1];
  assign T121 = T122 == 1'h1;
  assign T122 = io_inChannels_2_flit_x[1'h0:1'h0];
  assign T123 = T125 | T124;
  assign T124 = ~ io_inChannels_2_flitValid;
  assign T125 = T126 & T114;
  assign T126 = RouterBuffer_4_io_enq_ready & io_inChannels_2_flitValid;
  assign T128 = T129 | reset;
  assign T129 = T131 | T130;
  assign T130 = T1099 & T114;
  assign T131 = ~ T1099;
  assign T133 = T134 | reset;
  assign T134 = T145 | T135;
  assign T135 = ~ T136;
  assign T136 = T137 == 1'h1;
  assign T137 = T138;
  assign T138 = T143 ? T141 : T139;
  assign T139 = T140[6'h24:6'h24];
  assign T140 = io_inChannels_1_flit_x[6'h36:1'h1];
  assign T141 = T142[4'hd:4'hd];
  assign T142 = io_inChannels_1_flit_x[5'h1f:1'h1];
  assign T143 = T144 == 1'h1;
  assign T144 = io_inChannels_1_flit_x[1'h0:1'h0];
  assign T145 = T147 | T146;
  assign T146 = ~ io_inChannels_1_flitValid;
  assign T147 = T148 & T136;
  assign T148 = RouterBuffer_3_io_enq_ready & io_inChannels_1_flitValid;
  assign T150 = T151 | reset;
  assign T151 = T153 | T152;
  assign T152 = T1243 & T136;
  assign T153 = ~ T1243;
  assign T155 = T156 | reset;
  assign T156 = T167 | T157;
  assign T157 = ~ T158;
  assign T158 = T159 == 1'h0;
  assign T159 = T160;
  assign T160 = T165 ? T163 : T161;
  assign T161 = T162[6'h24:6'h24];
  assign T162 = io_inChannels_1_flit_x[6'h36:1'h1];
  assign T163 = T164[4'hd:4'hd];
  assign T164 = io_inChannels_1_flit_x[5'h1f:1'h1];
  assign T165 = T166 == 1'h1;
  assign T166 = io_inChannels_1_flit_x[1'h0:1'h0];
  assign T167 = T169 | T168;
  assign T168 = ~ io_inChannels_1_flitValid;
  assign T169 = T170 & T158;
  assign T170 = RouterBuffer_2_io_enq_ready & io_inChannels_1_flitValid;
  assign T172 = T173 | reset;
  assign T173 = T175 | T174;
  assign T174 = T1387 & T158;
  assign T175 = ~ T1387;
  assign T177 = T178 | reset;
  assign T178 = T189 | T179;
  assign T179 = ~ T180;
  assign T180 = T181 == 1'h1;
  assign T181 = T182;
  assign T182 = T187 ? T185 : T183;
  assign T183 = T184[6'h24:6'h24];
  assign T184 = io_inChannels_0_flit_x[6'h36:1'h1];
  assign T185 = T186[4'hd:4'hd];
  assign T186 = io_inChannels_0_flit_x[5'h1f:1'h1];
  assign T187 = T188 == 1'h1;
  assign T188 = io_inChannels_0_flit_x[1'h0:1'h0];
  assign T189 = T191 | T190;
  assign T190 = ~ io_inChannels_0_flitValid;
  assign T191 = T192 & T180;
  assign T192 = RouterBuffer_1_io_enq_ready & io_inChannels_0_flitValid;
  assign T194 = T195 | reset;
  assign T195 = T197 | T196;
  assign T196 = T1531 & T180;
  assign T197 = ~ T1531;
  assign T199 = T200 | reset;
  assign T200 = T211 | T201;
  assign T201 = ~ T202;
  assign T202 = T203 == 1'h0;
  assign T203 = T204;
  assign T204 = T209 ? T207 : T205;
  assign T205 = T206[6'h24:6'h24];
  assign T206 = io_inChannels_0_flit_x[6'h36:1'h1];
  assign T207 = T208[4'hd:4'hd];
  assign T208 = io_inChannels_0_flit_x[5'h1f:1'h1];
  assign T209 = T210 == 1'h1;
  assign T210 = io_inChannels_0_flit_x[1'h0:1'h0];
  assign T211 = T213 | T212;
  assign T212 = ~ io_inChannels_0_flitValid;
  assign T213 = T214 & T202;
  assign T214 = RouterBuffer_io_enq_ready & io_inChannels_0_flitValid;
  assign T216 = T217 | reset;
  assign T217 = T219 | T218;
  assign T218 = T1675 & T202;
  assign T219 = ~ T1675;
  assign T220 = T1722 & T221;
  assign T221 = T222 == 1'h1;
  assign T222 = T223;
  assign T223 = T228 ? T226 : T224;
  assign T224 = T225[6'h24:6'h24];
  assign T225 = switch_io_outPorts_4_x[6'h36:1'h1];
  assign T226 = T227[4'hd:4'hd];
  assign T227 = switch_io_outPorts_4_x[5'h1f:1'h1];
  assign T228 = T229 == 1'h1;
  assign T229 = switch_io_outPorts_4_x[1'h0:1'h0];
  assign T230 = T1722 & T231;
  assign T231 = T222 == 1'h0;
  assign T232 = T1905 & T233;
  assign T233 = T234 == 1'h1;
  assign T234 = T235;
  assign T235 = T240 ? T238 : T236;
  assign T236 = T237[6'h24:6'h24];
  assign T237 = switch_io_outPorts_3_x[6'h36:1'h1];
  assign T238 = T239[4'hd:4'hd];
  assign T239 = switch_io_outPorts_3_x[5'h1f:1'h1];
  assign T240 = T241 == 1'h1;
  assign T241 = switch_io_outPorts_3_x[1'h0:1'h0];
  assign T242 = T1905 & T243;
  assign T243 = T234 == 1'h0;
  assign T244 = T1968 & T245;
  assign T245 = T246 == 1'h1;
  assign T246 = T247;
  assign T247 = T252 ? T250 : T248;
  assign T248 = T249[6'h24:6'h24];
  assign T249 = switch_io_outPorts_2_x[6'h36:1'h1];
  assign T250 = T251[4'hd:4'hd];
  assign T251 = switch_io_outPorts_2_x[5'h1f:1'h1];
  assign T252 = T253 == 1'h1;
  assign T253 = switch_io_outPorts_2_x[1'h0:1'h0];
  assign T254 = T1968 & T255;
  assign T255 = T246 == 1'h0;
  assign T256 = T2031 & T257;
  assign T257 = T258 == 1'h1;
  assign T258 = T259;
  assign T259 = T264 ? T262 : T260;
  assign T260 = T261[6'h24:6'h24];
  assign T261 = switch_io_outPorts_1_x[6'h36:1'h1];
  assign T262 = T263[4'hd:4'hd];
  assign T263 = switch_io_outPorts_1_x[5'h1f:1'h1];
  assign T264 = T265 == 1'h1;
  assign T265 = switch_io_outPorts_1_x[1'h0:1'h0];
  assign T266 = T2031 & T267;
  assign T267 = T258 == 1'h0;
  assign T268 = T2094 & T269;
  assign T269 = T270 == 1'h1;
  assign T270 = T271;
  assign T271 = T276 ? T274 : T272;
  assign T272 = T273[6'h24:6'h24];
  assign T273 = switch_io_outPorts_0_x[6'h36:1'h1];
  assign T274 = T275[4'hd:4'hd];
  assign T275 = switch_io_outPorts_0_x[5'h1f:1'h1];
  assign T276 = T277 == 1'h1;
  assign T277 = switch_io_outPorts_0_x[1'h0:1'h0];
  assign T278 = T2094 & T279;
  assign T279 = T270 == 1'h0;
  assign T280 = T281;
  assign T281 = io_inChannels_4_flit_x;
  assign T3112 = R282[1'h0:1'h0];
  assign T3113 = reset ? 55'h0 : T283;
  assign T283 = T284 ? T3114 : R282;
  assign T3114 = {51'h0, vcAllocator_io_chosens_9};
  assign T284 = T285 & vcAllocator_io_resources_9_valid;
  assign T285 = VCRouterStateManagement_9_io_currentState == 3'h2;
  assign T286 = T287;
  assign T287 = RouterBuffer_9_io_deq_bits_x;
  assign T288 = T300 | T289;
  assign T289 = T290 == 2'h1;
  assign T290 = T299 ? VCRouterOutputStateManagement_4_io_currentState : T291;
  assign T291 = T298 ? T296 : T292;
  assign T292 = T293 ? VCRouterOutputStateManagement_1_io_currentState : VCRouterOutputStateManagement_io_currentState;
  assign T293 = T294[1'h0:1'h0];
  assign T294 = R295;
  assign T3115 = reset ? 3'h0 : CMeshDOR_9_io_result;
  assign T296 = T297 ? VCRouterOutputStateManagement_3_io_currentState : VCRouterOutputStateManagement_2_io_currentState;
  assign T297 = T294[1'h0:1'h0];
  assign T298 = T294[1'h1:1'h1];
  assign T299 = T294[2'h2:2'h2];
  assign T300 = T290 == 2'h2;
  assign T301 = T319 ? T311 : T302;
  assign T302 = T310 ? creditConsReady_4_0 : T303;
  assign T303 = T309 ? T307 : T304;
  assign T304 = T305 ? creditConsReady_1_0 : creditConsReady_0_0;
  assign creditConsReady_0_0 = CreditCon_io_outCredit;
  assign creditConsReady_1_0 = CreditCon_2_io_outCredit;
  assign T305 = T306[1'h0:1'h0];
  assign T306 = R295;
  assign T307 = T308 ? creditConsReady_3_0 : creditConsReady_2_0;
  assign creditConsReady_2_0 = CreditCon_4_io_outCredit;
  assign creditConsReady_3_0 = CreditCon_6_io_outCredit;
  assign T308 = T306[1'h0:1'h0];
  assign T309 = T306[1'h1:1'h1];
  assign creditConsReady_4_0 = CreditCon_8_io_outCredit;
  assign T310 = T306[2'h2:2'h2];
  assign T311 = T318 ? creditConsReady_4_1 : T312;
  assign T312 = T317 ? T315 : T313;
  assign T313 = T314 ? creditConsReady_1_1 : creditConsReady_0_1;
  assign creditConsReady_0_1 = CreditCon_1_io_outCredit;
  assign creditConsReady_1_1 = CreditCon_3_io_outCredit;
  assign T314 = T306[1'h0:1'h0];
  assign T315 = T316 ? creditConsReady_3_1 : creditConsReady_2_1;
  assign creditConsReady_2_1 = CreditCon_5_io_outCredit;
  assign creditConsReady_3_1 = CreditCon_7_io_outCredit;
  assign T316 = T306[1'h0:1'h0];
  assign T317 = T306[1'h1:1'h1];
  assign creditConsReady_4_1 = CreditCon_9_io_outCredit;
  assign T318 = T306[2'h2:2'h2];
  assign T319 = T3116;
  assign T3116 = R282[1'h0:1'h0];
  assign T320 = T331 & T321;
  assign T321 = T322 == 4'h9;
  assign T322 = T330 ? swAllocator_io_chosens_4 : T323;
  assign T323 = T329 ? T327 : T324;
  assign T324 = T325 ? swAllocator_io_chosens_1 : swAllocator_io_chosens_0;
  assign T325 = T326[1'h0:1'h0];
  assign T326 = R295;
  assign T327 = T328 ? swAllocator_io_chosens_3 : swAllocator_io_chosens_2;
  assign T328 = T326[1'h0:1'h0];
  assign T329 = T326[1'h1:1'h1];
  assign T330 = T326[2'h2:2'h2];
  assign T331 = T339 ? swAllocator_io_requests_4_9_grant : T332;
  assign T332 = T338 ? T336 : T333;
  assign T333 = T334 ? swAllocator_io_requests_1_9_grant : swAllocator_io_requests_0_9_grant;
  assign T334 = T335[1'h0:1'h0];
  assign T335 = R295;
  assign T336 = T337 ? swAllocator_io_requests_3_9_grant : swAllocator_io_requests_2_9_grant;
  assign T337 = T335[1'h0:1'h0];
  assign T338 = T335[1'h1:1'h1];
  assign T339 = T335[2'h2:2'h2];
  assign T340 = RouterBuffer_9_io_deq_valid & T341;
  assign T341 = T342;
  assign T342 = T347 ? T345 : T343;
  assign T343 = T344[6'h25:6'h25];
  assign T344 = RouterBuffer_9_io_deq_bits_x[6'h36:1'h1];
  assign T345 = T346[4'he:4'he];
  assign T346 = RouterBuffer_9_io_deq_bits_x[5'h1f:1'h1];
  assign T347 = T348 == 1'h1;
  assign T348 = RouterBuffer_9_io_deq_bits_x[1'h0:1'h0];
  assign T3117 = reset ? 1'h0 : RouterBuffer_9_io_deq_valid;
  assign T350 = T351[2'h2:1'h0];
  assign T351 = T352[5'h1f:1'h1];
  assign T352 = RouterRegFile_9_io_readData;
  assign T353 = T351[3'h4:2'h3];
  assign T354 = T351[3'h6:3'h5];
  assign T355 = T351[4'h8:3'h7];
  assign T356 = T351[4'hc:4'h9];
  assign T357 = T351[4'hd:4'hd];
  assign T358 = T351[4'he:4'he];
  assign T359 = T351[5'h1e:4'hf];
  assign T360 = T374 ? T371 : T361;
  assign T361 = T367 ? 1'h0 : T362;
  assign T362 = T363 & T301;
  assign T363 = T365 & T364;
  assign T364 = VCRouterStateManagement_9_io_currentState == 3'h4;
  assign T365 = T320 | T366;
  assign T366 = VCRouterStateManagement_9_io_currentState == 3'h4;
  assign T367 = T369 & T368;
  assign T368 = ~ RouterRegFile_9_io_readValid;
  assign T369 = T370 == 1'h1;
  assign T370 = RouterBuffer_9_io_deq_bits_x[1'h0:1'h0];
  assign T371 = T372 & T301;
  assign T372 = T365 & T373;
  assign T373 = 3'h3 <= VCRouterStateManagement_9_io_currentState;
  assign T374 = T378 & T375;
  assign T375 = T376 & RouterRegFile_9_io_readValid;
  assign T376 = T377 == 1'h1;
  assign T377 = RouterBuffer_9_io_deq_bits_x[1'h0:1'h0];
  assign T378 = T367 ^ 1'h1;
  assign T379 = io_inChannels_4_flitValid & T4;
  assign T380 = T381 & RouterRegFile_9_io_readValid;
  assign T381 = RouterRegFile_9_io_rvPipelineReg_0 ^ 1'h1;
  assign T382 = T384 & T383;
  assign T383 = VCRouterStateManagement_9_io_currentState == 3'h2;
  assign T384 = RouterRegFile_9_io_rvPipelineReg_0 & vcAllocator_io_resources_9_valid;
  assign T385 = T387 & T386;
  assign T386 = VCRouterStateManagement_9_io_currentState == 3'h3;
  assign T387 = RouterRegFile_9_io_rvPipelineReg_1 & T320;
  assign T3118 = {24'h0, T388};
  assign T388 = T389;
  assign T389 = {T393, T390};
  assign T390 = {T392, T391};
  assign T391 = {CMeshDOR_9_io_outHeadFlit_destination_0, CMeshDOR_9_io_outHeadFlit_priorityLevel};
  assign T392 = {CMeshDOR_9_io_outHeadFlit_destination_2, CMeshDOR_9_io_outHeadFlit_destination_1};
  assign T393 = {T395, T394};
  assign T394 = {CMeshDOR_9_io_outHeadFlit_vcPort, CMeshDOR_9_io_outHeadFlit_packetType};
  assign T395 = {CMeshDOR_9_io_outHeadFlit_packetID, CMeshDOR_9_io_outHeadFlit_isTail};
  assign T396 = T398 & T397;
  assign T397 = VCRouterStateManagement_9_io_currentState == 3'h4;
  assign T398 = T399 & T301;
  assign T399 = T365 & flitsAreTail_9;
  assign flitsAreTail_9 = T400;
  assign T400 = T401 & RouterBuffer_9_io_deq_valid;
  assign T401 = T402;
  assign T402 = T407 ? T405 : T403;
  assign T403 = T404[6'h25:6'h25];
  assign T404 = RouterBuffer_9_io_deq_bits_x[6'h36:1'h1];
  assign T405 = T406[4'he:4'he];
  assign T406 = RouterBuffer_9_io_deq_bits_x[5'h1f:1'h1];
  assign T407 = T408 == 1'h1;
  assign T408 = RouterBuffer_9_io_deq_bits_x[1'h0:1'h0];
  assign T409 = T410 ? T379 : 1'h0;
  assign T410 = T411 == 1'h1;
  assign T411 = io_inChannels_4_flit_x[1'h0:1'h0];
  assign T412 = T410 ? T413 : 55'h0;
  assign T413 = io_inChannels_4_flit_x;
  assign T414 = T374 ? T420 : T415;
  assign T415 = T367 ? 1'h0 : T416;
  assign T416 = T417 & RouterBuffer_9_io_deq_valid;
  assign T417 = T418 & T301;
  assign T418 = T365 & T419;
  assign T419 = VCRouterStateManagement_9_io_currentState == 3'h4;
  assign T420 = T421 & RouterBuffer_9_io_deq_valid;
  assign T421 = T422 & T301;
  assign T422 = T365 & T423;
  assign T423 = 3'h3 <= VCRouterStateManagement_9_io_currentState;
  assign T424 = T425;
  assign T425 = io_inChannels_4_flit_x;
  assign T3119 = R426[1'h0:1'h0];
  assign T3120 = reset ? 55'h0 : T427;
  assign T427 = T428 ? T3121 : R426;
  assign T3121 = {51'h0, vcAllocator_io_chosens_8};
  assign T428 = T429 & vcAllocator_io_resources_8_valid;
  assign T429 = VCRouterStateManagement_8_io_currentState == 3'h2;
  assign T430 = T431;
  assign T431 = RouterBuffer_8_io_deq_bits_x;
  assign T432 = T444 | T433;
  assign T433 = T434 == 2'h1;
  assign T434 = T443 ? VCRouterOutputStateManagement_4_io_currentState : T435;
  assign T435 = T442 ? T440 : T436;
  assign T436 = T437 ? VCRouterOutputStateManagement_1_io_currentState : VCRouterOutputStateManagement_io_currentState;
  assign T437 = T438[1'h0:1'h0];
  assign T438 = R439;
  assign T3122 = reset ? 3'h0 : CMeshDOR_8_io_result;
  assign T440 = T441 ? VCRouterOutputStateManagement_3_io_currentState : VCRouterOutputStateManagement_2_io_currentState;
  assign T441 = T438[1'h0:1'h0];
  assign T442 = T438[1'h1:1'h1];
  assign T443 = T438[2'h2:2'h2];
  assign T444 = T434 == 2'h2;
  assign T445 = T463 ? T455 : T446;
  assign T446 = T454 ? creditConsReady_4_0 : T447;
  assign T447 = T453 ? T451 : T448;
  assign T448 = T449 ? creditConsReady_1_0 : creditConsReady_0_0;
  assign T449 = T450[1'h0:1'h0];
  assign T450 = R439;
  assign T451 = T452 ? creditConsReady_3_0 : creditConsReady_2_0;
  assign T452 = T450[1'h0:1'h0];
  assign T453 = T450[1'h1:1'h1];
  assign T454 = T450[2'h2:2'h2];
  assign T455 = T462 ? creditConsReady_4_1 : T456;
  assign T456 = T461 ? T459 : T457;
  assign T457 = T458 ? creditConsReady_1_1 : creditConsReady_0_1;
  assign T458 = T450[1'h0:1'h0];
  assign T459 = T460 ? creditConsReady_3_1 : creditConsReady_2_1;
  assign T460 = T450[1'h0:1'h0];
  assign T461 = T450[1'h1:1'h1];
  assign T462 = T450[2'h2:2'h2];
  assign T463 = T3123;
  assign T3123 = R426[1'h0:1'h0];
  assign T464 = T475 & T465;
  assign T465 = T466 == 4'h8;
  assign T466 = T474 ? swAllocator_io_chosens_4 : T467;
  assign T467 = T473 ? T471 : T468;
  assign T468 = T469 ? swAllocator_io_chosens_1 : swAllocator_io_chosens_0;
  assign T469 = T470[1'h0:1'h0];
  assign T470 = R439;
  assign T471 = T472 ? swAllocator_io_chosens_3 : swAllocator_io_chosens_2;
  assign T472 = T470[1'h0:1'h0];
  assign T473 = T470[1'h1:1'h1];
  assign T474 = T470[2'h2:2'h2];
  assign T475 = T483 ? swAllocator_io_requests_4_8_grant : T476;
  assign T476 = T482 ? T480 : T477;
  assign T477 = T478 ? swAllocator_io_requests_1_8_grant : swAllocator_io_requests_0_8_grant;
  assign T478 = T479[1'h0:1'h0];
  assign T479 = R439;
  assign T480 = T481 ? swAllocator_io_requests_3_8_grant : swAllocator_io_requests_2_8_grant;
  assign T481 = T479[1'h0:1'h0];
  assign T482 = T479[1'h1:1'h1];
  assign T483 = T479[2'h2:2'h2];
  assign T484 = RouterBuffer_8_io_deq_valid & T485;
  assign T485 = T486;
  assign T486 = T491 ? T489 : T487;
  assign T487 = T488[6'h25:6'h25];
  assign T488 = RouterBuffer_8_io_deq_bits_x[6'h36:1'h1];
  assign T489 = T490[4'he:4'he];
  assign T490 = RouterBuffer_8_io_deq_bits_x[5'h1f:1'h1];
  assign T491 = T492 == 1'h1;
  assign T492 = RouterBuffer_8_io_deq_bits_x[1'h0:1'h0];
  assign T3124 = reset ? 1'h0 : RouterBuffer_8_io_deq_valid;
  assign T494 = T495[2'h2:1'h0];
  assign T495 = T496[5'h1f:1'h1];
  assign T496 = RouterRegFile_8_io_readData;
  assign T497 = T495[3'h4:2'h3];
  assign T498 = T495[3'h6:3'h5];
  assign T499 = T495[4'h8:3'h7];
  assign T500 = T495[4'hc:4'h9];
  assign T501 = T495[4'hd:4'hd];
  assign T502 = T495[4'he:4'he];
  assign T503 = T495[5'h1e:4'hf];
  assign T504 = T518 ? T515 : T505;
  assign T505 = T511 ? 1'h0 : T506;
  assign T506 = T507 & T445;
  assign T507 = T509 & T508;
  assign T508 = VCRouterStateManagement_8_io_currentState == 3'h4;
  assign T509 = T464 | T510;
  assign T510 = VCRouterStateManagement_8_io_currentState == 3'h4;
  assign T511 = T513 & T512;
  assign T512 = ~ RouterRegFile_8_io_readValid;
  assign T513 = T514 == 1'h1;
  assign T514 = RouterBuffer_8_io_deq_bits_x[1'h0:1'h0];
  assign T515 = T516 & T445;
  assign T516 = T509 & T517;
  assign T517 = 3'h3 <= VCRouterStateManagement_8_io_currentState;
  assign T518 = T522 & T519;
  assign T519 = T520 & RouterRegFile_8_io_readValid;
  assign T520 = T521 == 1'h1;
  assign T521 = RouterBuffer_8_io_deq_bits_x[1'h0:1'h0];
  assign T522 = T511 ^ 1'h1;
  assign T523 = io_inChannels_4_flitValid & T26;
  assign T524 = T525 & RouterRegFile_8_io_readValid;
  assign T525 = RouterRegFile_8_io_rvPipelineReg_0 ^ 1'h1;
  assign T526 = T528 & T527;
  assign T527 = VCRouterStateManagement_8_io_currentState == 3'h2;
  assign T528 = RouterRegFile_8_io_rvPipelineReg_0 & vcAllocator_io_resources_8_valid;
  assign T529 = T531 & T530;
  assign T530 = VCRouterStateManagement_8_io_currentState == 3'h3;
  assign T531 = RouterRegFile_8_io_rvPipelineReg_1 & T464;
  assign T3125 = {24'h0, T532};
  assign T532 = T533;
  assign T533 = {T537, T534};
  assign T534 = {T536, T535};
  assign T535 = {CMeshDOR_8_io_outHeadFlit_destination_0, CMeshDOR_8_io_outHeadFlit_priorityLevel};
  assign T536 = {CMeshDOR_8_io_outHeadFlit_destination_2, CMeshDOR_8_io_outHeadFlit_destination_1};
  assign T537 = {T539, T538};
  assign T538 = {CMeshDOR_8_io_outHeadFlit_vcPort, CMeshDOR_8_io_outHeadFlit_packetType};
  assign T539 = {CMeshDOR_8_io_outHeadFlit_packetID, CMeshDOR_8_io_outHeadFlit_isTail};
  assign T540 = T542 & T541;
  assign T541 = VCRouterStateManagement_8_io_currentState == 3'h4;
  assign T542 = T543 & T445;
  assign T543 = T509 & flitsAreTail_8;
  assign flitsAreTail_8 = T544;
  assign T544 = T545 & RouterBuffer_8_io_deq_valid;
  assign T545 = T546;
  assign T546 = T551 ? T549 : T547;
  assign T547 = T548[6'h25:6'h25];
  assign T548 = RouterBuffer_8_io_deq_bits_x[6'h36:1'h1];
  assign T549 = T550[4'he:4'he];
  assign T550 = RouterBuffer_8_io_deq_bits_x[5'h1f:1'h1];
  assign T551 = T552 == 1'h1;
  assign T552 = RouterBuffer_8_io_deq_bits_x[1'h0:1'h0];
  assign T553 = T554 ? T523 : 1'h0;
  assign T554 = T555 == 1'h1;
  assign T555 = io_inChannels_4_flit_x[1'h0:1'h0];
  assign T556 = T554 ? T557 : 55'h0;
  assign T557 = io_inChannels_4_flit_x;
  assign T558 = T518 ? T564 : T559;
  assign T559 = T511 ? 1'h0 : T560;
  assign T560 = T561 & RouterBuffer_8_io_deq_valid;
  assign T561 = T562 & T445;
  assign T562 = T509 & T563;
  assign T563 = VCRouterStateManagement_8_io_currentState == 3'h4;
  assign T564 = T565 & RouterBuffer_8_io_deq_valid;
  assign T565 = T566 & T445;
  assign T566 = T509 & T567;
  assign T567 = 3'h3 <= VCRouterStateManagement_8_io_currentState;
  assign T568 = T569;
  assign T569 = io_inChannels_3_flit_x;
  assign T3126 = R570[1'h0:1'h0];
  assign T3127 = reset ? 55'h0 : T571;
  assign T571 = T572 ? T3128 : R570;
  assign T3128 = {51'h0, vcAllocator_io_chosens_7};
  assign T572 = T573 & vcAllocator_io_resources_7_valid;
  assign T573 = VCRouterStateManagement_7_io_currentState == 3'h2;
  assign T574 = T575;
  assign T575 = RouterBuffer_7_io_deq_bits_x;
  assign T576 = T588 | T577;
  assign T577 = T578 == 2'h1;
  assign T578 = T587 ? VCRouterOutputStateManagement_4_io_currentState : T579;
  assign T579 = T586 ? T584 : T580;
  assign T580 = T581 ? VCRouterOutputStateManagement_1_io_currentState : VCRouterOutputStateManagement_io_currentState;
  assign T581 = T582[1'h0:1'h0];
  assign T582 = R583;
  assign T3129 = reset ? 3'h0 : CMeshDOR_7_io_result;
  assign T584 = T585 ? VCRouterOutputStateManagement_3_io_currentState : VCRouterOutputStateManagement_2_io_currentState;
  assign T585 = T582[1'h0:1'h0];
  assign T586 = T582[1'h1:1'h1];
  assign T587 = T582[2'h2:2'h2];
  assign T588 = T578 == 2'h2;
  assign T589 = T607 ? T599 : T590;
  assign T590 = T598 ? creditConsReady_4_0 : T591;
  assign T591 = T597 ? T595 : T592;
  assign T592 = T593 ? creditConsReady_1_0 : creditConsReady_0_0;
  assign T593 = T594[1'h0:1'h0];
  assign T594 = R583;
  assign T595 = T596 ? creditConsReady_3_0 : creditConsReady_2_0;
  assign T596 = T594[1'h0:1'h0];
  assign T597 = T594[1'h1:1'h1];
  assign T598 = T594[2'h2:2'h2];
  assign T599 = T606 ? creditConsReady_4_1 : T600;
  assign T600 = T605 ? T603 : T601;
  assign T601 = T602 ? creditConsReady_1_1 : creditConsReady_0_1;
  assign T602 = T594[1'h0:1'h0];
  assign T603 = T604 ? creditConsReady_3_1 : creditConsReady_2_1;
  assign T604 = T594[1'h0:1'h0];
  assign T605 = T594[1'h1:1'h1];
  assign T606 = T594[2'h2:2'h2];
  assign T607 = T3130;
  assign T3130 = R570[1'h0:1'h0];
  assign T608 = T619 & T609;
  assign T609 = T610 == 4'h7;
  assign T610 = T618 ? swAllocator_io_chosens_4 : T611;
  assign T611 = T617 ? T615 : T612;
  assign T612 = T613 ? swAllocator_io_chosens_1 : swAllocator_io_chosens_0;
  assign T613 = T614[1'h0:1'h0];
  assign T614 = R583;
  assign T615 = T616 ? swAllocator_io_chosens_3 : swAllocator_io_chosens_2;
  assign T616 = T614[1'h0:1'h0];
  assign T617 = T614[1'h1:1'h1];
  assign T618 = T614[2'h2:2'h2];
  assign T619 = T627 ? swAllocator_io_requests_4_7_grant : T620;
  assign T620 = T626 ? T624 : T621;
  assign T621 = T622 ? swAllocator_io_requests_1_7_grant : swAllocator_io_requests_0_7_grant;
  assign T622 = T623[1'h0:1'h0];
  assign T623 = R583;
  assign T624 = T625 ? swAllocator_io_requests_3_7_grant : swAllocator_io_requests_2_7_grant;
  assign T625 = T623[1'h0:1'h0];
  assign T626 = T623[1'h1:1'h1];
  assign T627 = T623[2'h2:2'h2];
  assign T628 = RouterBuffer_7_io_deq_valid & T629;
  assign T629 = T630;
  assign T630 = T635 ? T633 : T631;
  assign T631 = T632[6'h25:6'h25];
  assign T632 = RouterBuffer_7_io_deq_bits_x[6'h36:1'h1];
  assign T633 = T634[4'he:4'he];
  assign T634 = RouterBuffer_7_io_deq_bits_x[5'h1f:1'h1];
  assign T635 = T636 == 1'h1;
  assign T636 = RouterBuffer_7_io_deq_bits_x[1'h0:1'h0];
  assign T3131 = reset ? 1'h0 : RouterBuffer_7_io_deq_valid;
  assign T638 = T639[2'h2:1'h0];
  assign T639 = T640[5'h1f:1'h1];
  assign T640 = RouterRegFile_7_io_readData;
  assign T641 = T639[3'h4:2'h3];
  assign T642 = T639[3'h6:3'h5];
  assign T643 = T639[4'h8:3'h7];
  assign T644 = T639[4'hc:4'h9];
  assign T645 = T639[4'hd:4'hd];
  assign T646 = T639[4'he:4'he];
  assign T647 = T639[5'h1e:4'hf];
  assign T648 = T662 ? T659 : T649;
  assign T649 = T655 ? 1'h0 : T650;
  assign T650 = T651 & T589;
  assign T651 = T653 & T652;
  assign T652 = VCRouterStateManagement_7_io_currentState == 3'h4;
  assign T653 = T608 | T654;
  assign T654 = VCRouterStateManagement_7_io_currentState == 3'h4;
  assign T655 = T657 & T656;
  assign T656 = ~ RouterRegFile_7_io_readValid;
  assign T657 = T658 == 1'h1;
  assign T658 = RouterBuffer_7_io_deq_bits_x[1'h0:1'h0];
  assign T659 = T660 & T589;
  assign T660 = T653 & T661;
  assign T661 = 3'h3 <= VCRouterStateManagement_7_io_currentState;
  assign T662 = T666 & T663;
  assign T663 = T664 & RouterRegFile_7_io_readValid;
  assign T664 = T665 == 1'h1;
  assign T665 = RouterBuffer_7_io_deq_bits_x[1'h0:1'h0];
  assign T666 = T655 ^ 1'h1;
  assign T667 = io_inChannels_3_flitValid & T48;
  assign T668 = T669 & RouterRegFile_7_io_readValid;
  assign T669 = RouterRegFile_7_io_rvPipelineReg_0 ^ 1'h1;
  assign T670 = T672 & T671;
  assign T671 = VCRouterStateManagement_7_io_currentState == 3'h2;
  assign T672 = RouterRegFile_7_io_rvPipelineReg_0 & vcAllocator_io_resources_7_valid;
  assign T673 = T675 & T674;
  assign T674 = VCRouterStateManagement_7_io_currentState == 3'h3;
  assign T675 = RouterRegFile_7_io_rvPipelineReg_1 & T608;
  assign T3132 = {24'h0, T676};
  assign T676 = T677;
  assign T677 = {T681, T678};
  assign T678 = {T680, T679};
  assign T679 = {CMeshDOR_7_io_outHeadFlit_destination_0, CMeshDOR_7_io_outHeadFlit_priorityLevel};
  assign T680 = {CMeshDOR_7_io_outHeadFlit_destination_2, CMeshDOR_7_io_outHeadFlit_destination_1};
  assign T681 = {T683, T682};
  assign T682 = {CMeshDOR_7_io_outHeadFlit_vcPort, CMeshDOR_7_io_outHeadFlit_packetType};
  assign T683 = {CMeshDOR_7_io_outHeadFlit_packetID, CMeshDOR_7_io_outHeadFlit_isTail};
  assign T684 = T686 & T685;
  assign T685 = VCRouterStateManagement_7_io_currentState == 3'h4;
  assign T686 = T687 & T589;
  assign T687 = T653 & flitsAreTail_7;
  assign flitsAreTail_7 = T688;
  assign T688 = T689 & RouterBuffer_7_io_deq_valid;
  assign T689 = T690;
  assign T690 = T695 ? T693 : T691;
  assign T691 = T692[6'h25:6'h25];
  assign T692 = RouterBuffer_7_io_deq_bits_x[6'h36:1'h1];
  assign T693 = T694[4'he:4'he];
  assign T694 = RouterBuffer_7_io_deq_bits_x[5'h1f:1'h1];
  assign T695 = T696 == 1'h1;
  assign T696 = RouterBuffer_7_io_deq_bits_x[1'h0:1'h0];
  assign T697 = T698 ? T667 : 1'h0;
  assign T698 = T699 == 1'h1;
  assign T699 = io_inChannels_3_flit_x[1'h0:1'h0];
  assign T700 = T698 ? T701 : 55'h0;
  assign T701 = io_inChannels_3_flit_x;
  assign T702 = T662 ? T708 : T703;
  assign T703 = T655 ? 1'h0 : T704;
  assign T704 = T705 & RouterBuffer_7_io_deq_valid;
  assign T705 = T706 & T589;
  assign T706 = T653 & T707;
  assign T707 = VCRouterStateManagement_7_io_currentState == 3'h4;
  assign T708 = T709 & RouterBuffer_7_io_deq_valid;
  assign T709 = T710 & T589;
  assign T710 = T653 & T711;
  assign T711 = 3'h3 <= VCRouterStateManagement_7_io_currentState;
  assign T712 = T713;
  assign T713 = io_inChannels_3_flit_x;
  assign T3133 = R714[1'h0:1'h0];
  assign T3134 = reset ? 55'h0 : T715;
  assign T715 = T716 ? T3135 : R714;
  assign T3135 = {51'h0, vcAllocator_io_chosens_6};
  assign T716 = T717 & vcAllocator_io_resources_6_valid;
  assign T717 = VCRouterStateManagement_6_io_currentState == 3'h2;
  assign T718 = T719;
  assign T719 = RouterBuffer_6_io_deq_bits_x;
  assign T720 = T732 | T721;
  assign T721 = T722 == 2'h1;
  assign T722 = T731 ? VCRouterOutputStateManagement_4_io_currentState : T723;
  assign T723 = T730 ? T728 : T724;
  assign T724 = T725 ? VCRouterOutputStateManagement_1_io_currentState : VCRouterOutputStateManagement_io_currentState;
  assign T725 = T726[1'h0:1'h0];
  assign T726 = R727;
  assign T3136 = reset ? 3'h0 : CMeshDOR_6_io_result;
  assign T728 = T729 ? VCRouterOutputStateManagement_3_io_currentState : VCRouterOutputStateManagement_2_io_currentState;
  assign T729 = T726[1'h0:1'h0];
  assign T730 = T726[1'h1:1'h1];
  assign T731 = T726[2'h2:2'h2];
  assign T732 = T722 == 2'h2;
  assign T733 = T751 ? T743 : T734;
  assign T734 = T742 ? creditConsReady_4_0 : T735;
  assign T735 = T741 ? T739 : T736;
  assign T736 = T737 ? creditConsReady_1_0 : creditConsReady_0_0;
  assign T737 = T738[1'h0:1'h0];
  assign T738 = R727;
  assign T739 = T740 ? creditConsReady_3_0 : creditConsReady_2_0;
  assign T740 = T738[1'h0:1'h0];
  assign T741 = T738[1'h1:1'h1];
  assign T742 = T738[2'h2:2'h2];
  assign T743 = T750 ? creditConsReady_4_1 : T744;
  assign T744 = T749 ? T747 : T745;
  assign T745 = T746 ? creditConsReady_1_1 : creditConsReady_0_1;
  assign T746 = T738[1'h0:1'h0];
  assign T747 = T748 ? creditConsReady_3_1 : creditConsReady_2_1;
  assign T748 = T738[1'h0:1'h0];
  assign T749 = T738[1'h1:1'h1];
  assign T750 = T738[2'h2:2'h2];
  assign T751 = T3137;
  assign T3137 = R714[1'h0:1'h0];
  assign T752 = T763 & T753;
  assign T753 = T754 == 4'h6;
  assign T754 = T762 ? swAllocator_io_chosens_4 : T755;
  assign T755 = T761 ? T759 : T756;
  assign T756 = T757 ? swAllocator_io_chosens_1 : swAllocator_io_chosens_0;
  assign T757 = T758[1'h0:1'h0];
  assign T758 = R727;
  assign T759 = T760 ? swAllocator_io_chosens_3 : swAllocator_io_chosens_2;
  assign T760 = T758[1'h0:1'h0];
  assign T761 = T758[1'h1:1'h1];
  assign T762 = T758[2'h2:2'h2];
  assign T763 = T771 ? swAllocator_io_requests_4_6_grant : T764;
  assign T764 = T770 ? T768 : T765;
  assign T765 = T766 ? swAllocator_io_requests_1_6_grant : swAllocator_io_requests_0_6_grant;
  assign T766 = T767[1'h0:1'h0];
  assign T767 = R727;
  assign T768 = T769 ? swAllocator_io_requests_3_6_grant : swAllocator_io_requests_2_6_grant;
  assign T769 = T767[1'h0:1'h0];
  assign T770 = T767[1'h1:1'h1];
  assign T771 = T767[2'h2:2'h2];
  assign T772 = RouterBuffer_6_io_deq_valid & T773;
  assign T773 = T774;
  assign T774 = T779 ? T777 : T775;
  assign T775 = T776[6'h25:6'h25];
  assign T776 = RouterBuffer_6_io_deq_bits_x[6'h36:1'h1];
  assign T777 = T778[4'he:4'he];
  assign T778 = RouterBuffer_6_io_deq_bits_x[5'h1f:1'h1];
  assign T779 = T780 == 1'h1;
  assign T780 = RouterBuffer_6_io_deq_bits_x[1'h0:1'h0];
  assign T3138 = reset ? 1'h0 : RouterBuffer_6_io_deq_valid;
  assign T782 = T783[2'h2:1'h0];
  assign T783 = T784[5'h1f:1'h1];
  assign T784 = RouterRegFile_6_io_readData;
  assign T785 = T783[3'h4:2'h3];
  assign T786 = T783[3'h6:3'h5];
  assign T787 = T783[4'h8:3'h7];
  assign T788 = T783[4'hc:4'h9];
  assign T789 = T783[4'hd:4'hd];
  assign T790 = T783[4'he:4'he];
  assign T791 = T783[5'h1e:4'hf];
  assign T792 = T806 ? T803 : T793;
  assign T793 = T799 ? 1'h0 : T794;
  assign T794 = T795 & T733;
  assign T795 = T797 & T796;
  assign T796 = VCRouterStateManagement_6_io_currentState == 3'h4;
  assign T797 = T752 | T798;
  assign T798 = VCRouterStateManagement_6_io_currentState == 3'h4;
  assign T799 = T801 & T800;
  assign T800 = ~ RouterRegFile_6_io_readValid;
  assign T801 = T802 == 1'h1;
  assign T802 = RouterBuffer_6_io_deq_bits_x[1'h0:1'h0];
  assign T803 = T804 & T733;
  assign T804 = T797 & T805;
  assign T805 = 3'h3 <= VCRouterStateManagement_6_io_currentState;
  assign T806 = T810 & T807;
  assign T807 = T808 & RouterRegFile_6_io_readValid;
  assign T808 = T809 == 1'h1;
  assign T809 = RouterBuffer_6_io_deq_bits_x[1'h0:1'h0];
  assign T810 = T799 ^ 1'h1;
  assign T811 = io_inChannels_3_flitValid & T70;
  assign T812 = T813 & RouterRegFile_6_io_readValid;
  assign T813 = RouterRegFile_6_io_rvPipelineReg_0 ^ 1'h1;
  assign T814 = T816 & T815;
  assign T815 = VCRouterStateManagement_6_io_currentState == 3'h2;
  assign T816 = RouterRegFile_6_io_rvPipelineReg_0 & vcAllocator_io_resources_6_valid;
  assign T817 = T819 & T818;
  assign T818 = VCRouterStateManagement_6_io_currentState == 3'h3;
  assign T819 = RouterRegFile_6_io_rvPipelineReg_1 & T752;
  assign T3139 = {24'h0, T820};
  assign T820 = T821;
  assign T821 = {T825, T822};
  assign T822 = {T824, T823};
  assign T823 = {CMeshDOR_6_io_outHeadFlit_destination_0, CMeshDOR_6_io_outHeadFlit_priorityLevel};
  assign T824 = {CMeshDOR_6_io_outHeadFlit_destination_2, CMeshDOR_6_io_outHeadFlit_destination_1};
  assign T825 = {T827, T826};
  assign T826 = {CMeshDOR_6_io_outHeadFlit_vcPort, CMeshDOR_6_io_outHeadFlit_packetType};
  assign T827 = {CMeshDOR_6_io_outHeadFlit_packetID, CMeshDOR_6_io_outHeadFlit_isTail};
  assign T828 = T830 & T829;
  assign T829 = VCRouterStateManagement_6_io_currentState == 3'h4;
  assign T830 = T831 & T733;
  assign T831 = T797 & flitsAreTail_6;
  assign flitsAreTail_6 = T832;
  assign T832 = T833 & RouterBuffer_6_io_deq_valid;
  assign T833 = T834;
  assign T834 = T839 ? T837 : T835;
  assign T835 = T836[6'h25:6'h25];
  assign T836 = RouterBuffer_6_io_deq_bits_x[6'h36:1'h1];
  assign T837 = T838[4'he:4'he];
  assign T838 = RouterBuffer_6_io_deq_bits_x[5'h1f:1'h1];
  assign T839 = T840 == 1'h1;
  assign T840 = RouterBuffer_6_io_deq_bits_x[1'h0:1'h0];
  assign T841 = T842 ? T811 : 1'h0;
  assign T842 = T843 == 1'h1;
  assign T843 = io_inChannels_3_flit_x[1'h0:1'h0];
  assign T844 = T842 ? T845 : 55'h0;
  assign T845 = io_inChannels_3_flit_x;
  assign T846 = T806 ? T852 : T847;
  assign T847 = T799 ? 1'h0 : T848;
  assign T848 = T849 & RouterBuffer_6_io_deq_valid;
  assign T849 = T850 & T733;
  assign T850 = T797 & T851;
  assign T851 = VCRouterStateManagement_6_io_currentState == 3'h4;
  assign T852 = T853 & RouterBuffer_6_io_deq_valid;
  assign T853 = T854 & T733;
  assign T854 = T797 & T855;
  assign T855 = 3'h3 <= VCRouterStateManagement_6_io_currentState;
  assign T856 = T857;
  assign T857 = io_inChannels_2_flit_x;
  assign T3140 = R858[1'h0:1'h0];
  assign T3141 = reset ? 55'h0 : T859;
  assign T859 = T860 ? T3142 : R858;
  assign T3142 = {51'h0, vcAllocator_io_chosens_5};
  assign T860 = T861 & vcAllocator_io_resources_5_valid;
  assign T861 = VCRouterStateManagement_5_io_currentState == 3'h2;
  assign T862 = T863;
  assign T863 = RouterBuffer_5_io_deq_bits_x;
  assign T864 = T876 | T865;
  assign T865 = T866 == 2'h1;
  assign T866 = T875 ? VCRouterOutputStateManagement_4_io_currentState : T867;
  assign T867 = T874 ? T872 : T868;
  assign T868 = T869 ? VCRouterOutputStateManagement_1_io_currentState : VCRouterOutputStateManagement_io_currentState;
  assign T869 = T870[1'h0:1'h0];
  assign T870 = R871;
  assign T3143 = reset ? 3'h0 : CMeshDOR_5_io_result;
  assign T872 = T873 ? VCRouterOutputStateManagement_3_io_currentState : VCRouterOutputStateManagement_2_io_currentState;
  assign T873 = T870[1'h0:1'h0];
  assign T874 = T870[1'h1:1'h1];
  assign T875 = T870[2'h2:2'h2];
  assign T876 = T866 == 2'h2;
  assign T877 = T895 ? T887 : T878;
  assign T878 = T886 ? creditConsReady_4_0 : T879;
  assign T879 = T885 ? T883 : T880;
  assign T880 = T881 ? creditConsReady_1_0 : creditConsReady_0_0;
  assign T881 = T882[1'h0:1'h0];
  assign T882 = R871;
  assign T883 = T884 ? creditConsReady_3_0 : creditConsReady_2_0;
  assign T884 = T882[1'h0:1'h0];
  assign T885 = T882[1'h1:1'h1];
  assign T886 = T882[2'h2:2'h2];
  assign T887 = T894 ? creditConsReady_4_1 : T888;
  assign T888 = T893 ? T891 : T889;
  assign T889 = T890 ? creditConsReady_1_1 : creditConsReady_0_1;
  assign T890 = T882[1'h0:1'h0];
  assign T891 = T892 ? creditConsReady_3_1 : creditConsReady_2_1;
  assign T892 = T882[1'h0:1'h0];
  assign T893 = T882[1'h1:1'h1];
  assign T894 = T882[2'h2:2'h2];
  assign T895 = T3144;
  assign T3144 = R858[1'h0:1'h0];
  assign T896 = T907 & T897;
  assign T897 = T898 == 4'h5;
  assign T898 = T906 ? swAllocator_io_chosens_4 : T899;
  assign T899 = T905 ? T903 : T900;
  assign T900 = T901 ? swAllocator_io_chosens_1 : swAllocator_io_chosens_0;
  assign T901 = T902[1'h0:1'h0];
  assign T902 = R871;
  assign T903 = T904 ? swAllocator_io_chosens_3 : swAllocator_io_chosens_2;
  assign T904 = T902[1'h0:1'h0];
  assign T905 = T902[1'h1:1'h1];
  assign T906 = T902[2'h2:2'h2];
  assign T907 = T915 ? swAllocator_io_requests_4_5_grant : T908;
  assign T908 = T914 ? T912 : T909;
  assign T909 = T910 ? swAllocator_io_requests_1_5_grant : swAllocator_io_requests_0_5_grant;
  assign T910 = T911[1'h0:1'h0];
  assign T911 = R871;
  assign T912 = T913 ? swAllocator_io_requests_3_5_grant : swAllocator_io_requests_2_5_grant;
  assign T913 = T911[1'h0:1'h0];
  assign T914 = T911[1'h1:1'h1];
  assign T915 = T911[2'h2:2'h2];
  assign T916 = RouterBuffer_5_io_deq_valid & T917;
  assign T917 = T918;
  assign T918 = T923 ? T921 : T919;
  assign T919 = T920[6'h25:6'h25];
  assign T920 = RouterBuffer_5_io_deq_bits_x[6'h36:1'h1];
  assign T921 = T922[4'he:4'he];
  assign T922 = RouterBuffer_5_io_deq_bits_x[5'h1f:1'h1];
  assign T923 = T924 == 1'h1;
  assign T924 = RouterBuffer_5_io_deq_bits_x[1'h0:1'h0];
  assign T3145 = reset ? 1'h0 : RouterBuffer_5_io_deq_valid;
  assign T926 = T927[2'h2:1'h0];
  assign T927 = T928[5'h1f:1'h1];
  assign T928 = RouterRegFile_5_io_readData;
  assign T929 = T927[3'h4:2'h3];
  assign T930 = T927[3'h6:3'h5];
  assign T931 = T927[4'h8:3'h7];
  assign T932 = T927[4'hc:4'h9];
  assign T933 = T927[4'hd:4'hd];
  assign T934 = T927[4'he:4'he];
  assign T935 = T927[5'h1e:4'hf];
  assign T936 = T950 ? T947 : T937;
  assign T937 = T943 ? 1'h0 : T938;
  assign T938 = T939 & T877;
  assign T939 = T941 & T940;
  assign T940 = VCRouterStateManagement_5_io_currentState == 3'h4;
  assign T941 = T896 | T942;
  assign T942 = VCRouterStateManagement_5_io_currentState == 3'h4;
  assign T943 = T945 & T944;
  assign T944 = ~ RouterRegFile_5_io_readValid;
  assign T945 = T946 == 1'h1;
  assign T946 = RouterBuffer_5_io_deq_bits_x[1'h0:1'h0];
  assign T947 = T948 & T877;
  assign T948 = T941 & T949;
  assign T949 = 3'h3 <= VCRouterStateManagement_5_io_currentState;
  assign T950 = T954 & T951;
  assign T951 = T952 & RouterRegFile_5_io_readValid;
  assign T952 = T953 == 1'h1;
  assign T953 = RouterBuffer_5_io_deq_bits_x[1'h0:1'h0];
  assign T954 = T943 ^ 1'h1;
  assign T955 = io_inChannels_2_flitValid & T92;
  assign T956 = T957 & RouterRegFile_5_io_readValid;
  assign T957 = RouterRegFile_5_io_rvPipelineReg_0 ^ 1'h1;
  assign T958 = T960 & T959;
  assign T959 = VCRouterStateManagement_5_io_currentState == 3'h2;
  assign T960 = RouterRegFile_5_io_rvPipelineReg_0 & vcAllocator_io_resources_5_valid;
  assign T961 = T963 & T962;
  assign T962 = VCRouterStateManagement_5_io_currentState == 3'h3;
  assign T963 = RouterRegFile_5_io_rvPipelineReg_1 & T896;
  assign T3146 = {24'h0, T964};
  assign T964 = T965;
  assign T965 = {T969, T966};
  assign T966 = {T968, T967};
  assign T967 = {CMeshDOR_5_io_outHeadFlit_destination_0, CMeshDOR_5_io_outHeadFlit_priorityLevel};
  assign T968 = {CMeshDOR_5_io_outHeadFlit_destination_2, CMeshDOR_5_io_outHeadFlit_destination_1};
  assign T969 = {T971, T970};
  assign T970 = {CMeshDOR_5_io_outHeadFlit_vcPort, CMeshDOR_5_io_outHeadFlit_packetType};
  assign T971 = {CMeshDOR_5_io_outHeadFlit_packetID, CMeshDOR_5_io_outHeadFlit_isTail};
  assign T972 = T974 & T973;
  assign T973 = VCRouterStateManagement_5_io_currentState == 3'h4;
  assign T974 = T975 & T877;
  assign T975 = T941 & flitsAreTail_5;
  assign flitsAreTail_5 = T976;
  assign T976 = T977 & RouterBuffer_5_io_deq_valid;
  assign T977 = T978;
  assign T978 = T983 ? T981 : T979;
  assign T979 = T980[6'h25:6'h25];
  assign T980 = RouterBuffer_5_io_deq_bits_x[6'h36:1'h1];
  assign T981 = T982[4'he:4'he];
  assign T982 = RouterBuffer_5_io_deq_bits_x[5'h1f:1'h1];
  assign T983 = T984 == 1'h1;
  assign T984 = RouterBuffer_5_io_deq_bits_x[1'h0:1'h0];
  assign T985 = T986 ? T955 : 1'h0;
  assign T986 = T987 == 1'h1;
  assign T987 = io_inChannels_2_flit_x[1'h0:1'h0];
  assign T988 = T986 ? T989 : 55'h0;
  assign T989 = io_inChannels_2_flit_x;
  assign T990 = T950 ? T996 : T991;
  assign T991 = T943 ? 1'h0 : T992;
  assign T992 = T993 & RouterBuffer_5_io_deq_valid;
  assign T993 = T994 & T877;
  assign T994 = T941 & T995;
  assign T995 = VCRouterStateManagement_5_io_currentState == 3'h4;
  assign T996 = T997 & RouterBuffer_5_io_deq_valid;
  assign T997 = T998 & T877;
  assign T998 = T941 & T999;
  assign T999 = 3'h3 <= VCRouterStateManagement_5_io_currentState;
  assign T1000 = T1001;
  assign T1001 = io_inChannels_2_flit_x;
  assign T3147 = R1002[1'h0:1'h0];
  assign T3148 = reset ? 55'h0 : T1003;
  assign T1003 = T1004 ? T3149 : R1002;
  assign T3149 = {51'h0, vcAllocator_io_chosens_4};
  assign T1004 = T1005 & vcAllocator_io_resources_4_valid;
  assign T1005 = VCRouterStateManagement_4_io_currentState == 3'h2;
  assign T1006 = T1007;
  assign T1007 = RouterBuffer_4_io_deq_bits_x;
  assign T1008 = T1020 | T1009;
  assign T1009 = T1010 == 2'h1;
  assign T1010 = T1019 ? VCRouterOutputStateManagement_4_io_currentState : T1011;
  assign T1011 = T1018 ? T1016 : T1012;
  assign T1012 = T1013 ? VCRouterOutputStateManagement_1_io_currentState : VCRouterOutputStateManagement_io_currentState;
  assign T1013 = T1014[1'h0:1'h0];
  assign T1014 = R1015;
  assign T3150 = reset ? 3'h0 : CMeshDOR_4_io_result;
  assign T1016 = T1017 ? VCRouterOutputStateManagement_3_io_currentState : VCRouterOutputStateManagement_2_io_currentState;
  assign T1017 = T1014[1'h0:1'h0];
  assign T1018 = T1014[1'h1:1'h1];
  assign T1019 = T1014[2'h2:2'h2];
  assign T1020 = T1010 == 2'h2;
  assign T1021 = T1039 ? T1031 : T1022;
  assign T1022 = T1030 ? creditConsReady_4_0 : T1023;
  assign T1023 = T1029 ? T1027 : T1024;
  assign T1024 = T1025 ? creditConsReady_1_0 : creditConsReady_0_0;
  assign T1025 = T1026[1'h0:1'h0];
  assign T1026 = R1015;
  assign T1027 = T1028 ? creditConsReady_3_0 : creditConsReady_2_0;
  assign T1028 = T1026[1'h0:1'h0];
  assign T1029 = T1026[1'h1:1'h1];
  assign T1030 = T1026[2'h2:2'h2];
  assign T1031 = T1038 ? creditConsReady_4_1 : T1032;
  assign T1032 = T1037 ? T1035 : T1033;
  assign T1033 = T1034 ? creditConsReady_1_1 : creditConsReady_0_1;
  assign T1034 = T1026[1'h0:1'h0];
  assign T1035 = T1036 ? creditConsReady_3_1 : creditConsReady_2_1;
  assign T1036 = T1026[1'h0:1'h0];
  assign T1037 = T1026[1'h1:1'h1];
  assign T1038 = T1026[2'h2:2'h2];
  assign T1039 = T3151;
  assign T3151 = R1002[1'h0:1'h0];
  assign T1040 = T1051 & T1041;
  assign T1041 = T1042 == 4'h4;
  assign T1042 = T1050 ? swAllocator_io_chosens_4 : T1043;
  assign T1043 = T1049 ? T1047 : T1044;
  assign T1044 = T1045 ? swAllocator_io_chosens_1 : swAllocator_io_chosens_0;
  assign T1045 = T1046[1'h0:1'h0];
  assign T1046 = R1015;
  assign T1047 = T1048 ? swAllocator_io_chosens_3 : swAllocator_io_chosens_2;
  assign T1048 = T1046[1'h0:1'h0];
  assign T1049 = T1046[1'h1:1'h1];
  assign T1050 = T1046[2'h2:2'h2];
  assign T1051 = T1059 ? swAllocator_io_requests_4_4_grant : T1052;
  assign T1052 = T1058 ? T1056 : T1053;
  assign T1053 = T1054 ? swAllocator_io_requests_1_4_grant : swAllocator_io_requests_0_4_grant;
  assign T1054 = T1055[1'h0:1'h0];
  assign T1055 = R1015;
  assign T1056 = T1057 ? swAllocator_io_requests_3_4_grant : swAllocator_io_requests_2_4_grant;
  assign T1057 = T1055[1'h0:1'h0];
  assign T1058 = T1055[1'h1:1'h1];
  assign T1059 = T1055[2'h2:2'h2];
  assign T1060 = RouterBuffer_4_io_deq_valid & T1061;
  assign T1061 = T1062;
  assign T1062 = T1067 ? T1065 : T1063;
  assign T1063 = T1064[6'h25:6'h25];
  assign T1064 = RouterBuffer_4_io_deq_bits_x[6'h36:1'h1];
  assign T1065 = T1066[4'he:4'he];
  assign T1066 = RouterBuffer_4_io_deq_bits_x[5'h1f:1'h1];
  assign T1067 = T1068 == 1'h1;
  assign T1068 = RouterBuffer_4_io_deq_bits_x[1'h0:1'h0];
  assign T3152 = reset ? 1'h0 : RouterBuffer_4_io_deq_valid;
  assign T1070 = T1071[2'h2:1'h0];
  assign T1071 = T1072[5'h1f:1'h1];
  assign T1072 = RouterRegFile_4_io_readData;
  assign T1073 = T1071[3'h4:2'h3];
  assign T1074 = T1071[3'h6:3'h5];
  assign T1075 = T1071[4'h8:3'h7];
  assign T1076 = T1071[4'hc:4'h9];
  assign T1077 = T1071[4'hd:4'hd];
  assign T1078 = T1071[4'he:4'he];
  assign T1079 = T1071[5'h1e:4'hf];
  assign T1080 = T1094 ? T1091 : T1081;
  assign T1081 = T1087 ? 1'h0 : T1082;
  assign T1082 = T1083 & T1021;
  assign T1083 = T1085 & T1084;
  assign T1084 = VCRouterStateManagement_4_io_currentState == 3'h4;
  assign T1085 = T1040 | T1086;
  assign T1086 = VCRouterStateManagement_4_io_currentState == 3'h4;
  assign T1087 = T1089 & T1088;
  assign T1088 = ~ RouterRegFile_4_io_readValid;
  assign T1089 = T1090 == 1'h1;
  assign T1090 = RouterBuffer_4_io_deq_bits_x[1'h0:1'h0];
  assign T1091 = T1092 & T1021;
  assign T1092 = T1085 & T1093;
  assign T1093 = 3'h3 <= VCRouterStateManagement_4_io_currentState;
  assign T1094 = T1098 & T1095;
  assign T1095 = T1096 & RouterRegFile_4_io_readValid;
  assign T1096 = T1097 == 1'h1;
  assign T1097 = RouterBuffer_4_io_deq_bits_x[1'h0:1'h0];
  assign T1098 = T1087 ^ 1'h1;
  assign T1099 = io_inChannels_2_flitValid & T114;
  assign T1100 = T1101 & RouterRegFile_4_io_readValid;
  assign T1101 = RouterRegFile_4_io_rvPipelineReg_0 ^ 1'h1;
  assign T1102 = T1104 & T1103;
  assign T1103 = VCRouterStateManagement_4_io_currentState == 3'h2;
  assign T1104 = RouterRegFile_4_io_rvPipelineReg_0 & vcAllocator_io_resources_4_valid;
  assign T1105 = T1107 & T1106;
  assign T1106 = VCRouterStateManagement_4_io_currentState == 3'h3;
  assign T1107 = RouterRegFile_4_io_rvPipelineReg_1 & T1040;
  assign T3153 = {24'h0, T1108};
  assign T1108 = T1109;
  assign T1109 = {T1113, T1110};
  assign T1110 = {T1112, T1111};
  assign T1111 = {CMeshDOR_4_io_outHeadFlit_destination_0, CMeshDOR_4_io_outHeadFlit_priorityLevel};
  assign T1112 = {CMeshDOR_4_io_outHeadFlit_destination_2, CMeshDOR_4_io_outHeadFlit_destination_1};
  assign T1113 = {T1115, T1114};
  assign T1114 = {CMeshDOR_4_io_outHeadFlit_vcPort, CMeshDOR_4_io_outHeadFlit_packetType};
  assign T1115 = {CMeshDOR_4_io_outHeadFlit_packetID, CMeshDOR_4_io_outHeadFlit_isTail};
  assign T1116 = T1118 & T1117;
  assign T1117 = VCRouterStateManagement_4_io_currentState == 3'h4;
  assign T1118 = T1119 & T1021;
  assign T1119 = T1085 & flitsAreTail_4;
  assign flitsAreTail_4 = T1120;
  assign T1120 = T1121 & RouterBuffer_4_io_deq_valid;
  assign T1121 = T1122;
  assign T1122 = T1127 ? T1125 : T1123;
  assign T1123 = T1124[6'h25:6'h25];
  assign T1124 = RouterBuffer_4_io_deq_bits_x[6'h36:1'h1];
  assign T1125 = T1126[4'he:4'he];
  assign T1126 = RouterBuffer_4_io_deq_bits_x[5'h1f:1'h1];
  assign T1127 = T1128 == 1'h1;
  assign T1128 = RouterBuffer_4_io_deq_bits_x[1'h0:1'h0];
  assign T1129 = T1130 ? T1099 : 1'h0;
  assign T1130 = T1131 == 1'h1;
  assign T1131 = io_inChannels_2_flit_x[1'h0:1'h0];
  assign T1132 = T1130 ? T1133 : 55'h0;
  assign T1133 = io_inChannels_2_flit_x;
  assign T1134 = T1094 ? T1140 : T1135;
  assign T1135 = T1087 ? 1'h0 : T1136;
  assign T1136 = T1137 & RouterBuffer_4_io_deq_valid;
  assign T1137 = T1138 & T1021;
  assign T1138 = T1085 & T1139;
  assign T1139 = VCRouterStateManagement_4_io_currentState == 3'h4;
  assign T1140 = T1141 & RouterBuffer_4_io_deq_valid;
  assign T1141 = T1142 & T1021;
  assign T1142 = T1085 & T1143;
  assign T1143 = 3'h3 <= VCRouterStateManagement_4_io_currentState;
  assign T1144 = T1145;
  assign T1145 = io_inChannels_1_flit_x;
  assign T3154 = R1146[1'h0:1'h0];
  assign T3155 = reset ? 55'h0 : T1147;
  assign T1147 = T1148 ? T3156 : R1146;
  assign T3156 = {51'h0, vcAllocator_io_chosens_3};
  assign T1148 = T1149 & vcAllocator_io_resources_3_valid;
  assign T1149 = VCRouterStateManagement_3_io_currentState == 3'h2;
  assign T1150 = T1151;
  assign T1151 = RouterBuffer_3_io_deq_bits_x;
  assign T1152 = T1164 | T1153;
  assign T1153 = T1154 == 2'h1;
  assign T1154 = T1163 ? VCRouterOutputStateManagement_4_io_currentState : T1155;
  assign T1155 = T1162 ? T1160 : T1156;
  assign T1156 = T1157 ? VCRouterOutputStateManagement_1_io_currentState : VCRouterOutputStateManagement_io_currentState;
  assign T1157 = T1158[1'h0:1'h0];
  assign T1158 = R1159;
  assign T3157 = reset ? 3'h0 : CMeshDOR_3_io_result;
  assign T1160 = T1161 ? VCRouterOutputStateManagement_3_io_currentState : VCRouterOutputStateManagement_2_io_currentState;
  assign T1161 = T1158[1'h0:1'h0];
  assign T1162 = T1158[1'h1:1'h1];
  assign T1163 = T1158[2'h2:2'h2];
  assign T1164 = T1154 == 2'h2;
  assign T1165 = T1183 ? T1175 : T1166;
  assign T1166 = T1174 ? creditConsReady_4_0 : T1167;
  assign T1167 = T1173 ? T1171 : T1168;
  assign T1168 = T1169 ? creditConsReady_1_0 : creditConsReady_0_0;
  assign T1169 = T1170[1'h0:1'h0];
  assign T1170 = R1159;
  assign T1171 = T1172 ? creditConsReady_3_0 : creditConsReady_2_0;
  assign T1172 = T1170[1'h0:1'h0];
  assign T1173 = T1170[1'h1:1'h1];
  assign T1174 = T1170[2'h2:2'h2];
  assign T1175 = T1182 ? creditConsReady_4_1 : T1176;
  assign T1176 = T1181 ? T1179 : T1177;
  assign T1177 = T1178 ? creditConsReady_1_1 : creditConsReady_0_1;
  assign T1178 = T1170[1'h0:1'h0];
  assign T1179 = T1180 ? creditConsReady_3_1 : creditConsReady_2_1;
  assign T1180 = T1170[1'h0:1'h0];
  assign T1181 = T1170[1'h1:1'h1];
  assign T1182 = T1170[2'h2:2'h2];
  assign T1183 = T3158;
  assign T3158 = R1146[1'h0:1'h0];
  assign T1184 = T1195 & T1185;
  assign T1185 = T1186 == 4'h3;
  assign T1186 = T1194 ? swAllocator_io_chosens_4 : T1187;
  assign T1187 = T1193 ? T1191 : T1188;
  assign T1188 = T1189 ? swAllocator_io_chosens_1 : swAllocator_io_chosens_0;
  assign T1189 = T1190[1'h0:1'h0];
  assign T1190 = R1159;
  assign T1191 = T1192 ? swAllocator_io_chosens_3 : swAllocator_io_chosens_2;
  assign T1192 = T1190[1'h0:1'h0];
  assign T1193 = T1190[1'h1:1'h1];
  assign T1194 = T1190[2'h2:2'h2];
  assign T1195 = T1203 ? swAllocator_io_requests_4_3_grant : T1196;
  assign T1196 = T1202 ? T1200 : T1197;
  assign T1197 = T1198 ? swAllocator_io_requests_1_3_grant : swAllocator_io_requests_0_3_grant;
  assign T1198 = T1199[1'h0:1'h0];
  assign T1199 = R1159;
  assign T1200 = T1201 ? swAllocator_io_requests_3_3_grant : swAllocator_io_requests_2_3_grant;
  assign T1201 = T1199[1'h0:1'h0];
  assign T1202 = T1199[1'h1:1'h1];
  assign T1203 = T1199[2'h2:2'h2];
  assign T1204 = RouterBuffer_3_io_deq_valid & T1205;
  assign T1205 = T1206;
  assign T1206 = T1211 ? T1209 : T1207;
  assign T1207 = T1208[6'h25:6'h25];
  assign T1208 = RouterBuffer_3_io_deq_bits_x[6'h36:1'h1];
  assign T1209 = T1210[4'he:4'he];
  assign T1210 = RouterBuffer_3_io_deq_bits_x[5'h1f:1'h1];
  assign T1211 = T1212 == 1'h1;
  assign T1212 = RouterBuffer_3_io_deq_bits_x[1'h0:1'h0];
  assign T3159 = reset ? 1'h0 : RouterBuffer_3_io_deq_valid;
  assign T1214 = T1215[2'h2:1'h0];
  assign T1215 = T1216[5'h1f:1'h1];
  assign T1216 = RouterRegFile_3_io_readData;
  assign T1217 = T1215[3'h4:2'h3];
  assign T1218 = T1215[3'h6:3'h5];
  assign T1219 = T1215[4'h8:3'h7];
  assign T1220 = T1215[4'hc:4'h9];
  assign T1221 = T1215[4'hd:4'hd];
  assign T1222 = T1215[4'he:4'he];
  assign T1223 = T1215[5'h1e:4'hf];
  assign T1224 = T1238 ? T1235 : T1225;
  assign T1225 = T1231 ? 1'h0 : T1226;
  assign T1226 = T1227 & T1165;
  assign T1227 = T1229 & T1228;
  assign T1228 = VCRouterStateManagement_3_io_currentState == 3'h4;
  assign T1229 = T1184 | T1230;
  assign T1230 = VCRouterStateManagement_3_io_currentState == 3'h4;
  assign T1231 = T1233 & T1232;
  assign T1232 = ~ RouterRegFile_3_io_readValid;
  assign T1233 = T1234 == 1'h1;
  assign T1234 = RouterBuffer_3_io_deq_bits_x[1'h0:1'h0];
  assign T1235 = T1236 & T1165;
  assign T1236 = T1229 & T1237;
  assign T1237 = 3'h3 <= VCRouterStateManagement_3_io_currentState;
  assign T1238 = T1242 & T1239;
  assign T1239 = T1240 & RouterRegFile_3_io_readValid;
  assign T1240 = T1241 == 1'h1;
  assign T1241 = RouterBuffer_3_io_deq_bits_x[1'h0:1'h0];
  assign T1242 = T1231 ^ 1'h1;
  assign T1243 = io_inChannels_1_flitValid & T136;
  assign T1244 = T1245 & RouterRegFile_3_io_readValid;
  assign T1245 = RouterRegFile_3_io_rvPipelineReg_0 ^ 1'h1;
  assign T1246 = T1248 & T1247;
  assign T1247 = VCRouterStateManagement_3_io_currentState == 3'h2;
  assign T1248 = RouterRegFile_3_io_rvPipelineReg_0 & vcAllocator_io_resources_3_valid;
  assign T1249 = T1251 & T1250;
  assign T1250 = VCRouterStateManagement_3_io_currentState == 3'h3;
  assign T1251 = RouterRegFile_3_io_rvPipelineReg_1 & T1184;
  assign T3160 = {24'h0, T1252};
  assign T1252 = T1253;
  assign T1253 = {T1257, T1254};
  assign T1254 = {T1256, T1255};
  assign T1255 = {CMeshDOR_3_io_outHeadFlit_destination_0, CMeshDOR_3_io_outHeadFlit_priorityLevel};
  assign T1256 = {CMeshDOR_3_io_outHeadFlit_destination_2, CMeshDOR_3_io_outHeadFlit_destination_1};
  assign T1257 = {T1259, T1258};
  assign T1258 = {CMeshDOR_3_io_outHeadFlit_vcPort, CMeshDOR_3_io_outHeadFlit_packetType};
  assign T1259 = {CMeshDOR_3_io_outHeadFlit_packetID, CMeshDOR_3_io_outHeadFlit_isTail};
  assign T1260 = T1262 & T1261;
  assign T1261 = VCRouterStateManagement_3_io_currentState == 3'h4;
  assign T1262 = T1263 & T1165;
  assign T1263 = T1229 & flitsAreTail_3;
  assign flitsAreTail_3 = T1264;
  assign T1264 = T1265 & RouterBuffer_3_io_deq_valid;
  assign T1265 = T1266;
  assign T1266 = T1271 ? T1269 : T1267;
  assign T1267 = T1268[6'h25:6'h25];
  assign T1268 = RouterBuffer_3_io_deq_bits_x[6'h36:1'h1];
  assign T1269 = T1270[4'he:4'he];
  assign T1270 = RouterBuffer_3_io_deq_bits_x[5'h1f:1'h1];
  assign T1271 = T1272 == 1'h1;
  assign T1272 = RouterBuffer_3_io_deq_bits_x[1'h0:1'h0];
  assign T1273 = T1274 ? T1243 : 1'h0;
  assign T1274 = T1275 == 1'h1;
  assign T1275 = io_inChannels_1_flit_x[1'h0:1'h0];
  assign T1276 = T1274 ? T1277 : 55'h0;
  assign T1277 = io_inChannels_1_flit_x;
  assign T1278 = T1238 ? T1284 : T1279;
  assign T1279 = T1231 ? 1'h0 : T1280;
  assign T1280 = T1281 & RouterBuffer_3_io_deq_valid;
  assign T1281 = T1282 & T1165;
  assign T1282 = T1229 & T1283;
  assign T1283 = VCRouterStateManagement_3_io_currentState == 3'h4;
  assign T1284 = T1285 & RouterBuffer_3_io_deq_valid;
  assign T1285 = T1286 & T1165;
  assign T1286 = T1229 & T1287;
  assign T1287 = 3'h3 <= VCRouterStateManagement_3_io_currentState;
  assign T1288 = T1289;
  assign T1289 = io_inChannels_1_flit_x;
  assign T3161 = R1290[1'h0:1'h0];
  assign T3162 = reset ? 55'h0 : T1291;
  assign T1291 = T1292 ? T3163 : R1290;
  assign T3163 = {51'h0, vcAllocator_io_chosens_2};
  assign T1292 = T1293 & vcAllocator_io_resources_2_valid;
  assign T1293 = VCRouterStateManagement_2_io_currentState == 3'h2;
  assign T1294 = T1295;
  assign T1295 = RouterBuffer_2_io_deq_bits_x;
  assign T1296 = T1308 | T1297;
  assign T1297 = T1298 == 2'h1;
  assign T1298 = T1307 ? VCRouterOutputStateManagement_4_io_currentState : T1299;
  assign T1299 = T1306 ? T1304 : T1300;
  assign T1300 = T1301 ? VCRouterOutputStateManagement_1_io_currentState : VCRouterOutputStateManagement_io_currentState;
  assign T1301 = T1302[1'h0:1'h0];
  assign T1302 = R1303;
  assign T3164 = reset ? 3'h0 : CMeshDOR_2_io_result;
  assign T1304 = T1305 ? VCRouterOutputStateManagement_3_io_currentState : VCRouterOutputStateManagement_2_io_currentState;
  assign T1305 = T1302[1'h0:1'h0];
  assign T1306 = T1302[1'h1:1'h1];
  assign T1307 = T1302[2'h2:2'h2];
  assign T1308 = T1298 == 2'h2;
  assign T1309 = T1327 ? T1319 : T1310;
  assign T1310 = T1318 ? creditConsReady_4_0 : T1311;
  assign T1311 = T1317 ? T1315 : T1312;
  assign T1312 = T1313 ? creditConsReady_1_0 : creditConsReady_0_0;
  assign T1313 = T1314[1'h0:1'h0];
  assign T1314 = R1303;
  assign T1315 = T1316 ? creditConsReady_3_0 : creditConsReady_2_0;
  assign T1316 = T1314[1'h0:1'h0];
  assign T1317 = T1314[1'h1:1'h1];
  assign T1318 = T1314[2'h2:2'h2];
  assign T1319 = T1326 ? creditConsReady_4_1 : T1320;
  assign T1320 = T1325 ? T1323 : T1321;
  assign T1321 = T1322 ? creditConsReady_1_1 : creditConsReady_0_1;
  assign T1322 = T1314[1'h0:1'h0];
  assign T1323 = T1324 ? creditConsReady_3_1 : creditConsReady_2_1;
  assign T1324 = T1314[1'h0:1'h0];
  assign T1325 = T1314[1'h1:1'h1];
  assign T1326 = T1314[2'h2:2'h2];
  assign T1327 = T3165;
  assign T3165 = R1290[1'h0:1'h0];
  assign T1328 = T1339 & T1329;
  assign T1329 = T1330 == 4'h2;
  assign T1330 = T1338 ? swAllocator_io_chosens_4 : T1331;
  assign T1331 = T1337 ? T1335 : T1332;
  assign T1332 = T1333 ? swAllocator_io_chosens_1 : swAllocator_io_chosens_0;
  assign T1333 = T1334[1'h0:1'h0];
  assign T1334 = R1303;
  assign T1335 = T1336 ? swAllocator_io_chosens_3 : swAllocator_io_chosens_2;
  assign T1336 = T1334[1'h0:1'h0];
  assign T1337 = T1334[1'h1:1'h1];
  assign T1338 = T1334[2'h2:2'h2];
  assign T1339 = T1347 ? swAllocator_io_requests_4_2_grant : T1340;
  assign T1340 = T1346 ? T1344 : T1341;
  assign T1341 = T1342 ? swAllocator_io_requests_1_2_grant : swAllocator_io_requests_0_2_grant;
  assign T1342 = T1343[1'h0:1'h0];
  assign T1343 = R1303;
  assign T1344 = T1345 ? swAllocator_io_requests_3_2_grant : swAllocator_io_requests_2_2_grant;
  assign T1345 = T1343[1'h0:1'h0];
  assign T1346 = T1343[1'h1:1'h1];
  assign T1347 = T1343[2'h2:2'h2];
  assign T1348 = RouterBuffer_2_io_deq_valid & T1349;
  assign T1349 = T1350;
  assign T1350 = T1355 ? T1353 : T1351;
  assign T1351 = T1352[6'h25:6'h25];
  assign T1352 = RouterBuffer_2_io_deq_bits_x[6'h36:1'h1];
  assign T1353 = T1354[4'he:4'he];
  assign T1354 = RouterBuffer_2_io_deq_bits_x[5'h1f:1'h1];
  assign T1355 = T1356 == 1'h1;
  assign T1356 = RouterBuffer_2_io_deq_bits_x[1'h0:1'h0];
  assign T3166 = reset ? 1'h0 : RouterBuffer_2_io_deq_valid;
  assign T1358 = T1359[2'h2:1'h0];
  assign T1359 = T1360[5'h1f:1'h1];
  assign T1360 = RouterRegFile_2_io_readData;
  assign T1361 = T1359[3'h4:2'h3];
  assign T1362 = T1359[3'h6:3'h5];
  assign T1363 = T1359[4'h8:3'h7];
  assign T1364 = T1359[4'hc:4'h9];
  assign T1365 = T1359[4'hd:4'hd];
  assign T1366 = T1359[4'he:4'he];
  assign T1367 = T1359[5'h1e:4'hf];
  assign T1368 = T1382 ? T1379 : T1369;
  assign T1369 = T1375 ? 1'h0 : T1370;
  assign T1370 = T1371 & T1309;
  assign T1371 = T1373 & T1372;
  assign T1372 = VCRouterStateManagement_2_io_currentState == 3'h4;
  assign T1373 = T1328 | T1374;
  assign T1374 = VCRouterStateManagement_2_io_currentState == 3'h4;
  assign T1375 = T1377 & T1376;
  assign T1376 = ~ RouterRegFile_2_io_readValid;
  assign T1377 = T1378 == 1'h1;
  assign T1378 = RouterBuffer_2_io_deq_bits_x[1'h0:1'h0];
  assign T1379 = T1380 & T1309;
  assign T1380 = T1373 & T1381;
  assign T1381 = 3'h3 <= VCRouterStateManagement_2_io_currentState;
  assign T1382 = T1386 & T1383;
  assign T1383 = T1384 & RouterRegFile_2_io_readValid;
  assign T1384 = T1385 == 1'h1;
  assign T1385 = RouterBuffer_2_io_deq_bits_x[1'h0:1'h0];
  assign T1386 = T1375 ^ 1'h1;
  assign T1387 = io_inChannels_1_flitValid & T158;
  assign T1388 = T1389 & RouterRegFile_2_io_readValid;
  assign T1389 = RouterRegFile_2_io_rvPipelineReg_0 ^ 1'h1;
  assign T1390 = T1392 & T1391;
  assign T1391 = VCRouterStateManagement_2_io_currentState == 3'h2;
  assign T1392 = RouterRegFile_2_io_rvPipelineReg_0 & vcAllocator_io_resources_2_valid;
  assign T1393 = T1395 & T1394;
  assign T1394 = VCRouterStateManagement_2_io_currentState == 3'h3;
  assign T1395 = RouterRegFile_2_io_rvPipelineReg_1 & T1328;
  assign T3167 = {24'h0, T1396};
  assign T1396 = T1397;
  assign T1397 = {T1401, T1398};
  assign T1398 = {T1400, T1399};
  assign T1399 = {CMeshDOR_2_io_outHeadFlit_destination_0, CMeshDOR_2_io_outHeadFlit_priorityLevel};
  assign T1400 = {CMeshDOR_2_io_outHeadFlit_destination_2, CMeshDOR_2_io_outHeadFlit_destination_1};
  assign T1401 = {T1403, T1402};
  assign T1402 = {CMeshDOR_2_io_outHeadFlit_vcPort, CMeshDOR_2_io_outHeadFlit_packetType};
  assign T1403 = {CMeshDOR_2_io_outHeadFlit_packetID, CMeshDOR_2_io_outHeadFlit_isTail};
  assign T1404 = T1406 & T1405;
  assign T1405 = VCRouterStateManagement_2_io_currentState == 3'h4;
  assign T1406 = T1407 & T1309;
  assign T1407 = T1373 & flitsAreTail_2;
  assign flitsAreTail_2 = T1408;
  assign T1408 = T1409 & RouterBuffer_2_io_deq_valid;
  assign T1409 = T1410;
  assign T1410 = T1415 ? T1413 : T1411;
  assign T1411 = T1412[6'h25:6'h25];
  assign T1412 = RouterBuffer_2_io_deq_bits_x[6'h36:1'h1];
  assign T1413 = T1414[4'he:4'he];
  assign T1414 = RouterBuffer_2_io_deq_bits_x[5'h1f:1'h1];
  assign T1415 = T1416 == 1'h1;
  assign T1416 = RouterBuffer_2_io_deq_bits_x[1'h0:1'h0];
  assign T1417 = T1418 ? T1387 : 1'h0;
  assign T1418 = T1419 == 1'h1;
  assign T1419 = io_inChannels_1_flit_x[1'h0:1'h0];
  assign T1420 = T1418 ? T1421 : 55'h0;
  assign T1421 = io_inChannels_1_flit_x;
  assign T1422 = T1382 ? T1428 : T1423;
  assign T1423 = T1375 ? 1'h0 : T1424;
  assign T1424 = T1425 & RouterBuffer_2_io_deq_valid;
  assign T1425 = T1426 & T1309;
  assign T1426 = T1373 & T1427;
  assign T1427 = VCRouterStateManagement_2_io_currentState == 3'h4;
  assign T1428 = T1429 & RouterBuffer_2_io_deq_valid;
  assign T1429 = T1430 & T1309;
  assign T1430 = T1373 & T1431;
  assign T1431 = 3'h3 <= VCRouterStateManagement_2_io_currentState;
  assign T1432 = T1433;
  assign T1433 = io_inChannels_0_flit_x;
  assign T3168 = R1434[1'h0:1'h0];
  assign T3169 = reset ? 55'h0 : T1435;
  assign T1435 = T1436 ? T3170 : R1434;
  assign T3170 = {51'h0, vcAllocator_io_chosens_1};
  assign T1436 = T1437 & vcAllocator_io_resources_1_valid;
  assign T1437 = VCRouterStateManagement_1_io_currentState == 3'h2;
  assign T1438 = T1439;
  assign T1439 = RouterBuffer_1_io_deq_bits_x;
  assign T1440 = T1452 | T1441;
  assign T1441 = T1442 == 2'h1;
  assign T1442 = T1451 ? VCRouterOutputStateManagement_4_io_currentState : T1443;
  assign T1443 = T1450 ? T1448 : T1444;
  assign T1444 = T1445 ? VCRouterOutputStateManagement_1_io_currentState : VCRouterOutputStateManagement_io_currentState;
  assign T1445 = T1446[1'h0:1'h0];
  assign T1446 = R1447;
  assign T3171 = reset ? 3'h0 : CMeshDOR_1_io_result;
  assign T1448 = T1449 ? VCRouterOutputStateManagement_3_io_currentState : VCRouterOutputStateManagement_2_io_currentState;
  assign T1449 = T1446[1'h0:1'h0];
  assign T1450 = T1446[1'h1:1'h1];
  assign T1451 = T1446[2'h2:2'h2];
  assign T1452 = T1442 == 2'h2;
  assign T1453 = T1471 ? T1463 : T1454;
  assign T1454 = T1462 ? creditConsReady_4_0 : T1455;
  assign T1455 = T1461 ? T1459 : T1456;
  assign T1456 = T1457 ? creditConsReady_1_0 : creditConsReady_0_0;
  assign T1457 = T1458[1'h0:1'h0];
  assign T1458 = R1447;
  assign T1459 = T1460 ? creditConsReady_3_0 : creditConsReady_2_0;
  assign T1460 = T1458[1'h0:1'h0];
  assign T1461 = T1458[1'h1:1'h1];
  assign T1462 = T1458[2'h2:2'h2];
  assign T1463 = T1470 ? creditConsReady_4_1 : T1464;
  assign T1464 = T1469 ? T1467 : T1465;
  assign T1465 = T1466 ? creditConsReady_1_1 : creditConsReady_0_1;
  assign T1466 = T1458[1'h0:1'h0];
  assign T1467 = T1468 ? creditConsReady_3_1 : creditConsReady_2_1;
  assign T1468 = T1458[1'h0:1'h0];
  assign T1469 = T1458[1'h1:1'h1];
  assign T1470 = T1458[2'h2:2'h2];
  assign T1471 = T3172;
  assign T3172 = R1434[1'h0:1'h0];
  assign T1472 = T1483 & T1473;
  assign T1473 = T1474 == 4'h1;
  assign T1474 = T1482 ? swAllocator_io_chosens_4 : T1475;
  assign T1475 = T1481 ? T1479 : T1476;
  assign T1476 = T1477 ? swAllocator_io_chosens_1 : swAllocator_io_chosens_0;
  assign T1477 = T1478[1'h0:1'h0];
  assign T1478 = R1447;
  assign T1479 = T1480 ? swAllocator_io_chosens_3 : swAllocator_io_chosens_2;
  assign T1480 = T1478[1'h0:1'h0];
  assign T1481 = T1478[1'h1:1'h1];
  assign T1482 = T1478[2'h2:2'h2];
  assign T1483 = T1491 ? swAllocator_io_requests_4_1_grant : T1484;
  assign T1484 = T1490 ? T1488 : T1485;
  assign T1485 = T1486 ? swAllocator_io_requests_1_1_grant : swAllocator_io_requests_0_1_grant;
  assign T1486 = T1487[1'h0:1'h0];
  assign T1487 = R1447;
  assign T1488 = T1489 ? swAllocator_io_requests_3_1_grant : swAllocator_io_requests_2_1_grant;
  assign T1489 = T1487[1'h0:1'h0];
  assign T1490 = T1487[1'h1:1'h1];
  assign T1491 = T1487[2'h2:2'h2];
  assign T1492 = RouterBuffer_1_io_deq_valid & T1493;
  assign T1493 = T1494;
  assign T1494 = T1499 ? T1497 : T1495;
  assign T1495 = T1496[6'h25:6'h25];
  assign T1496 = RouterBuffer_1_io_deq_bits_x[6'h36:1'h1];
  assign T1497 = T1498[4'he:4'he];
  assign T1498 = RouterBuffer_1_io_deq_bits_x[5'h1f:1'h1];
  assign T1499 = T1500 == 1'h1;
  assign T1500 = RouterBuffer_1_io_deq_bits_x[1'h0:1'h0];
  assign T3173 = reset ? 1'h0 : RouterBuffer_1_io_deq_valid;
  assign T1502 = T1503[2'h2:1'h0];
  assign T1503 = T1504[5'h1f:1'h1];
  assign T1504 = RouterRegFile_1_io_readData;
  assign T1505 = T1503[3'h4:2'h3];
  assign T1506 = T1503[3'h6:3'h5];
  assign T1507 = T1503[4'h8:3'h7];
  assign T1508 = T1503[4'hc:4'h9];
  assign T1509 = T1503[4'hd:4'hd];
  assign T1510 = T1503[4'he:4'he];
  assign T1511 = T1503[5'h1e:4'hf];
  assign T1512 = T1526 ? T1523 : T1513;
  assign T1513 = T1519 ? 1'h0 : T1514;
  assign T1514 = T1515 & T1453;
  assign T1515 = T1517 & T1516;
  assign T1516 = VCRouterStateManagement_1_io_currentState == 3'h4;
  assign T1517 = T1472 | T1518;
  assign T1518 = VCRouterStateManagement_1_io_currentState == 3'h4;
  assign T1519 = T1521 & T1520;
  assign T1520 = ~ RouterRegFile_1_io_readValid;
  assign T1521 = T1522 == 1'h1;
  assign T1522 = RouterBuffer_1_io_deq_bits_x[1'h0:1'h0];
  assign T1523 = T1524 & T1453;
  assign T1524 = T1517 & T1525;
  assign T1525 = 3'h3 <= VCRouterStateManagement_1_io_currentState;
  assign T1526 = T1530 & T1527;
  assign T1527 = T1528 & RouterRegFile_1_io_readValid;
  assign T1528 = T1529 == 1'h1;
  assign T1529 = RouterBuffer_1_io_deq_bits_x[1'h0:1'h0];
  assign T1530 = T1519 ^ 1'h1;
  assign T1531 = io_inChannels_0_flitValid & T180;
  assign T1532 = T1533 & RouterRegFile_1_io_readValid;
  assign T1533 = RouterRegFile_1_io_rvPipelineReg_0 ^ 1'h1;
  assign T1534 = T1536 & T1535;
  assign T1535 = VCRouterStateManagement_1_io_currentState == 3'h2;
  assign T1536 = RouterRegFile_1_io_rvPipelineReg_0 & vcAllocator_io_resources_1_valid;
  assign T1537 = T1539 & T1538;
  assign T1538 = VCRouterStateManagement_1_io_currentState == 3'h3;
  assign T1539 = RouterRegFile_1_io_rvPipelineReg_1 & T1472;
  assign T3174 = {24'h0, T1540};
  assign T1540 = T1541;
  assign T1541 = {T1545, T1542};
  assign T1542 = {T1544, T1543};
  assign T1543 = {CMeshDOR_1_io_outHeadFlit_destination_0, CMeshDOR_1_io_outHeadFlit_priorityLevel};
  assign T1544 = {CMeshDOR_1_io_outHeadFlit_destination_2, CMeshDOR_1_io_outHeadFlit_destination_1};
  assign T1545 = {T1547, T1546};
  assign T1546 = {CMeshDOR_1_io_outHeadFlit_vcPort, CMeshDOR_1_io_outHeadFlit_packetType};
  assign T1547 = {CMeshDOR_1_io_outHeadFlit_packetID, CMeshDOR_1_io_outHeadFlit_isTail};
  assign T1548 = T1550 & T1549;
  assign T1549 = VCRouterStateManagement_1_io_currentState == 3'h4;
  assign T1550 = T1551 & T1453;
  assign T1551 = T1517 & flitsAreTail_1;
  assign flitsAreTail_1 = T1552;
  assign T1552 = T1553 & RouterBuffer_1_io_deq_valid;
  assign T1553 = T1554;
  assign T1554 = T1559 ? T1557 : T1555;
  assign T1555 = T1556[6'h25:6'h25];
  assign T1556 = RouterBuffer_1_io_deq_bits_x[6'h36:1'h1];
  assign T1557 = T1558[4'he:4'he];
  assign T1558 = RouterBuffer_1_io_deq_bits_x[5'h1f:1'h1];
  assign T1559 = T1560 == 1'h1;
  assign T1560 = RouterBuffer_1_io_deq_bits_x[1'h0:1'h0];
  assign T1561 = T1562 ? T1531 : 1'h0;
  assign T1562 = T1563 == 1'h1;
  assign T1563 = io_inChannels_0_flit_x[1'h0:1'h0];
  assign T1564 = T1562 ? T1565 : 55'h0;
  assign T1565 = io_inChannels_0_flit_x;
  assign T1566 = T1526 ? T1572 : T1567;
  assign T1567 = T1519 ? 1'h0 : T1568;
  assign T1568 = T1569 & RouterBuffer_1_io_deq_valid;
  assign T1569 = T1570 & T1453;
  assign T1570 = T1517 & T1571;
  assign T1571 = VCRouterStateManagement_1_io_currentState == 3'h4;
  assign T1572 = T1573 & RouterBuffer_1_io_deq_valid;
  assign T1573 = T1574 & T1453;
  assign T1574 = T1517 & T1575;
  assign T1575 = 3'h3 <= VCRouterStateManagement_1_io_currentState;
  assign T1576 = T1577;
  assign T1577 = io_inChannels_0_flit_x;
  assign T3175 = R1578[1'h0:1'h0];
  assign T3176 = reset ? 55'h0 : T1579;
  assign T1579 = T1580 ? T3177 : R1578;
  assign T3177 = {51'h0, vcAllocator_io_chosens_0};
  assign T1580 = T1581 & vcAllocator_io_resources_0_valid;
  assign T1581 = VCRouterStateManagement_io_currentState == 3'h2;
  assign T1582 = T1583;
  assign T1583 = RouterBuffer_io_deq_bits_x;
  assign T1584 = T1596 | T1585;
  assign T1585 = T1586 == 2'h1;
  assign T1586 = T1595 ? VCRouterOutputStateManagement_4_io_currentState : T1587;
  assign T1587 = T1594 ? T1592 : T1588;
  assign T1588 = T1589 ? VCRouterOutputStateManagement_1_io_currentState : VCRouterOutputStateManagement_io_currentState;
  assign T1589 = T1590[1'h0:1'h0];
  assign T1590 = R1591;
  assign T3178 = reset ? 3'h0 : CMeshDOR_io_result;
  assign T1592 = T1593 ? VCRouterOutputStateManagement_3_io_currentState : VCRouterOutputStateManagement_2_io_currentState;
  assign T1593 = T1590[1'h0:1'h0];
  assign T1594 = T1590[1'h1:1'h1];
  assign T1595 = T1590[2'h2:2'h2];
  assign T1596 = T1586 == 2'h2;
  assign T1597 = T1615 ? T1607 : T1598;
  assign T1598 = T1606 ? creditConsReady_4_0 : T1599;
  assign T1599 = T1605 ? T1603 : T1600;
  assign T1600 = T1601 ? creditConsReady_1_0 : creditConsReady_0_0;
  assign T1601 = T1602[1'h0:1'h0];
  assign T1602 = R1591;
  assign T1603 = T1604 ? creditConsReady_3_0 : creditConsReady_2_0;
  assign T1604 = T1602[1'h0:1'h0];
  assign T1605 = T1602[1'h1:1'h1];
  assign T1606 = T1602[2'h2:2'h2];
  assign T1607 = T1614 ? creditConsReady_4_1 : T1608;
  assign T1608 = T1613 ? T1611 : T1609;
  assign T1609 = T1610 ? creditConsReady_1_1 : creditConsReady_0_1;
  assign T1610 = T1602[1'h0:1'h0];
  assign T1611 = T1612 ? creditConsReady_3_1 : creditConsReady_2_1;
  assign T1612 = T1602[1'h0:1'h0];
  assign T1613 = T1602[1'h1:1'h1];
  assign T1614 = T1602[2'h2:2'h2];
  assign T1615 = T3179;
  assign T3179 = R1578[1'h0:1'h0];
  assign T1616 = T1627 & T1617;
  assign T1617 = T1618 == 4'h0;
  assign T1618 = T1626 ? swAllocator_io_chosens_4 : T1619;
  assign T1619 = T1625 ? T1623 : T1620;
  assign T1620 = T1621 ? swAllocator_io_chosens_1 : swAllocator_io_chosens_0;
  assign T1621 = T1622[1'h0:1'h0];
  assign T1622 = R1591;
  assign T1623 = T1624 ? swAllocator_io_chosens_3 : swAllocator_io_chosens_2;
  assign T1624 = T1622[1'h0:1'h0];
  assign T1625 = T1622[1'h1:1'h1];
  assign T1626 = T1622[2'h2:2'h2];
  assign T1627 = T1635 ? swAllocator_io_requests_4_0_grant : T1628;
  assign T1628 = T1634 ? T1632 : T1629;
  assign T1629 = T1630 ? swAllocator_io_requests_1_0_grant : swAllocator_io_requests_0_0_grant;
  assign T1630 = T1631[1'h0:1'h0];
  assign T1631 = R1591;
  assign T1632 = T1633 ? swAllocator_io_requests_3_0_grant : swAllocator_io_requests_2_0_grant;
  assign T1633 = T1631[1'h0:1'h0];
  assign T1634 = T1631[1'h1:1'h1];
  assign T1635 = T1631[2'h2:2'h2];
  assign T1636 = RouterBuffer_io_deq_valid & T1637;
  assign T1637 = T1638;
  assign T1638 = T1643 ? T1641 : T1639;
  assign T1639 = T1640[6'h25:6'h25];
  assign T1640 = RouterBuffer_io_deq_bits_x[6'h36:1'h1];
  assign T1641 = T1642[4'he:4'he];
  assign T1642 = RouterBuffer_io_deq_bits_x[5'h1f:1'h1];
  assign T1643 = T1644 == 1'h1;
  assign T1644 = RouterBuffer_io_deq_bits_x[1'h0:1'h0];
  assign T3180 = reset ? 1'h0 : RouterBuffer_io_deq_valid;
  assign T1646 = T1647[2'h2:1'h0];
  assign T1647 = T1648[5'h1f:1'h1];
  assign T1648 = RouterRegFile_io_readData;
  assign T1649 = T1647[3'h4:2'h3];
  assign T1650 = T1647[3'h6:3'h5];
  assign T1651 = T1647[4'h8:3'h7];
  assign T1652 = T1647[4'hc:4'h9];
  assign T1653 = T1647[4'hd:4'hd];
  assign T1654 = T1647[4'he:4'he];
  assign T1655 = T1647[5'h1e:4'hf];
  assign T1656 = T1670 ? T1667 : T1657;
  assign T1657 = T1663 ? 1'h0 : T1658;
  assign T1658 = T1659 & T1597;
  assign T1659 = T1661 & T1660;
  assign T1660 = VCRouterStateManagement_io_currentState == 3'h4;
  assign T1661 = T1616 | T1662;
  assign T1662 = VCRouterStateManagement_io_currentState == 3'h4;
  assign T1663 = T1665 & T1664;
  assign T1664 = ~ RouterRegFile_io_readValid;
  assign T1665 = T1666 == 1'h1;
  assign T1666 = RouterBuffer_io_deq_bits_x[1'h0:1'h0];
  assign T1667 = T1668 & T1597;
  assign T1668 = T1661 & T1669;
  assign T1669 = 3'h3 <= VCRouterStateManagement_io_currentState;
  assign T1670 = T1674 & T1671;
  assign T1671 = T1672 & RouterRegFile_io_readValid;
  assign T1672 = T1673 == 1'h1;
  assign T1673 = RouterBuffer_io_deq_bits_x[1'h0:1'h0];
  assign T1674 = T1663 ^ 1'h1;
  assign T1675 = io_inChannels_0_flitValid & T202;
  assign T1676 = T1677 & RouterRegFile_io_readValid;
  assign T1677 = RouterRegFile_io_rvPipelineReg_0 ^ 1'h1;
  assign T1678 = T1680 & T1679;
  assign T1679 = VCRouterStateManagement_io_currentState == 3'h2;
  assign T1680 = RouterRegFile_io_rvPipelineReg_0 & vcAllocator_io_resources_0_valid;
  assign T1681 = T1683 & T1682;
  assign T1682 = VCRouterStateManagement_io_currentState == 3'h3;
  assign T1683 = RouterRegFile_io_rvPipelineReg_1 & T1616;
  assign T3181 = {24'h0, T1684};
  assign T1684 = T1685;
  assign T1685 = {T1689, T1686};
  assign T1686 = {T1688, T1687};
  assign T1687 = {CMeshDOR_io_outHeadFlit_destination_0, CMeshDOR_io_outHeadFlit_priorityLevel};
  assign T1688 = {CMeshDOR_io_outHeadFlit_destination_2, CMeshDOR_io_outHeadFlit_destination_1};
  assign T1689 = {T1691, T1690};
  assign T1690 = {CMeshDOR_io_outHeadFlit_vcPort, CMeshDOR_io_outHeadFlit_packetType};
  assign T1691 = {CMeshDOR_io_outHeadFlit_packetID, CMeshDOR_io_outHeadFlit_isTail};
  assign T1692 = T1694 & T1693;
  assign T1693 = VCRouterStateManagement_io_currentState == 3'h4;
  assign T1694 = T1695 & T1597;
  assign T1695 = T1661 & flitsAreTail_0;
  assign flitsAreTail_0 = T1696;
  assign T1696 = T1697 & RouterBuffer_io_deq_valid;
  assign T1697 = T1698;
  assign T1698 = T1703 ? T1701 : T1699;
  assign T1699 = T1700[6'h25:6'h25];
  assign T1700 = RouterBuffer_io_deq_bits_x[6'h36:1'h1];
  assign T1701 = T1702[4'he:4'he];
  assign T1702 = RouterBuffer_io_deq_bits_x[5'h1f:1'h1];
  assign T1703 = T1704 == 1'h1;
  assign T1704 = RouterBuffer_io_deq_bits_x[1'h0:1'h0];
  assign T1705 = T1706 ? T1675 : 1'h0;
  assign T1706 = T1707 == 1'h1;
  assign T1707 = io_inChannels_0_flit_x[1'h0:1'h0];
  assign T1708 = T1706 ? T1709 : 55'h0;
  assign T1709 = io_inChannels_0_flit_x;
  assign T1710 = T1670 ? T1716 : T1711;
  assign T1711 = T1663 ? 1'h0 : T1712;
  assign T1712 = T1713 & RouterBuffer_io_deq_valid;
  assign T1713 = T1714 & T1597;
  assign T1714 = T1661 & T1715;
  assign T1715 = VCRouterStateManagement_io_currentState == 3'h4;
  assign T1716 = T1717 & RouterBuffer_io_deq_valid;
  assign T1717 = T1718 & T1597;
  assign T1718 = T1661 & T1719;
  assign T1719 = 3'h3 <= VCRouterStateManagement_io_currentState;
  assign T1720 = T1721 ? CreditCon_9_io_outCredit : CreditCon_8_io_outCredit;
  assign T1721 = T222;
  assign T1722 = T1723 != 10'h0;
  assign T1723 = T1724;
  assign T1724 = {T1814, T1725};
  assign T1725 = {T1779, T1726};
  assign T1726 = {readyToXmit_2_4, T1727};
  assign T1727 = {readyToXmit_1_4, readyToXmit_0_4};
  assign readyToXmit_0_4 = T1728;
  assign T1728 = T1742 ? T1738 : T1729;
  assign T1729 = T1734 ? T1730 : 1'h0;
  assign T1730 = T1731 & RouterBuffer_io_deq_valid;
  assign T1731 = T1732 & T1597;
  assign T1732 = T1661 & T1733;
  assign T1733 = 3'h3 <= VCRouterStateManagement_io_currentState;
  assign T1734 = T1670 & T1735;
  assign T1735 = T1736[3'h4:3'h4];
  assign T1736 = 1'h1 << T1737;
  assign T1737 = R1591;
  assign T1738 = T1739 & RouterBuffer_io_deq_valid;
  assign T1739 = T1740 & T1597;
  assign T1740 = T1661 & T1741;
  assign T1741 = VCRouterStateManagement_io_currentState == 3'h4;
  assign T1742 = T1743 & T1735;
  assign T1743 = T1744 ^ 1'h1;
  assign T1744 = T1663 | T1671;
  assign readyToXmit_1_4 = T1745;
  assign T1745 = T1759 ? T1755 : T1746;
  assign T1746 = T1751 ? T1747 : 1'h0;
  assign T1747 = T1748 & RouterBuffer_1_io_deq_valid;
  assign T1748 = T1749 & T1453;
  assign T1749 = T1517 & T1750;
  assign T1750 = 3'h3 <= VCRouterStateManagement_1_io_currentState;
  assign T1751 = T1526 & T1752;
  assign T1752 = T1753[3'h4:3'h4];
  assign T1753 = 1'h1 << T1754;
  assign T1754 = R1447;
  assign T1755 = T1756 & RouterBuffer_1_io_deq_valid;
  assign T1756 = T1757 & T1453;
  assign T1757 = T1517 & T1758;
  assign T1758 = VCRouterStateManagement_1_io_currentState == 3'h4;
  assign T1759 = T1760 & T1752;
  assign T1760 = T1761 ^ 1'h1;
  assign T1761 = T1519 | T1527;
  assign readyToXmit_2_4 = T1762;
  assign T1762 = T1776 ? T1772 : T1763;
  assign T1763 = T1768 ? T1764 : 1'h0;
  assign T1764 = T1765 & RouterBuffer_2_io_deq_valid;
  assign T1765 = T1766 & T1309;
  assign T1766 = T1373 & T1767;
  assign T1767 = 3'h3 <= VCRouterStateManagement_2_io_currentState;
  assign T1768 = T1382 & T1769;
  assign T1769 = T1770[3'h4:3'h4];
  assign T1770 = 1'h1 << T1771;
  assign T1771 = R1303;
  assign T1772 = T1773 & RouterBuffer_2_io_deq_valid;
  assign T1773 = T1774 & T1309;
  assign T1774 = T1373 & T1775;
  assign T1775 = VCRouterStateManagement_2_io_currentState == 3'h4;
  assign T1776 = T1777 & T1769;
  assign T1777 = T1778 ^ 1'h1;
  assign T1778 = T1375 | T1383;
  assign T1779 = {readyToXmit_4_4, readyToXmit_3_4};
  assign readyToXmit_3_4 = T1780;
  assign T1780 = T1794 ? T1790 : T1781;
  assign T1781 = T1786 ? T1782 : 1'h0;
  assign T1782 = T1783 & RouterBuffer_3_io_deq_valid;
  assign T1783 = T1784 & T1165;
  assign T1784 = T1229 & T1785;
  assign T1785 = 3'h3 <= VCRouterStateManagement_3_io_currentState;
  assign T1786 = T1238 & T1787;
  assign T1787 = T1788[3'h4:3'h4];
  assign T1788 = 1'h1 << T1789;
  assign T1789 = R1159;
  assign T1790 = T1791 & RouterBuffer_3_io_deq_valid;
  assign T1791 = T1792 & T1165;
  assign T1792 = T1229 & T1793;
  assign T1793 = VCRouterStateManagement_3_io_currentState == 3'h4;
  assign T1794 = T1795 & T1787;
  assign T1795 = T1796 ^ 1'h1;
  assign T1796 = T1231 | T1239;
  assign readyToXmit_4_4 = T1797;
  assign T1797 = T1811 ? T1807 : T1798;
  assign T1798 = T1803 ? T1799 : 1'h0;
  assign T1799 = T1800 & RouterBuffer_4_io_deq_valid;
  assign T1800 = T1801 & T1021;
  assign T1801 = T1085 & T1802;
  assign T1802 = 3'h3 <= VCRouterStateManagement_4_io_currentState;
  assign T1803 = T1094 & T1804;
  assign T1804 = T1805[3'h4:3'h4];
  assign T1805 = 1'h1 << T1806;
  assign T1806 = R1015;
  assign T1807 = T1808 & RouterBuffer_4_io_deq_valid;
  assign T1808 = T1809 & T1021;
  assign T1809 = T1085 & T1810;
  assign T1810 = VCRouterStateManagement_4_io_currentState == 3'h4;
  assign T1811 = T1812 & T1804;
  assign T1812 = T1813 ^ 1'h1;
  assign T1813 = T1087 | T1095;
  assign T1814 = {T1868, T1815};
  assign T1815 = {readyToXmit_7_4, T1816};
  assign T1816 = {readyToXmit_6_4, readyToXmit_5_4};
  assign readyToXmit_5_4 = T1817;
  assign T1817 = T1831 ? T1827 : T1818;
  assign T1818 = T1823 ? T1819 : 1'h0;
  assign T1819 = T1820 & RouterBuffer_5_io_deq_valid;
  assign T1820 = T1821 & T877;
  assign T1821 = T941 & T1822;
  assign T1822 = 3'h3 <= VCRouterStateManagement_5_io_currentState;
  assign T1823 = T950 & T1824;
  assign T1824 = T1825[3'h4:3'h4];
  assign T1825 = 1'h1 << T1826;
  assign T1826 = R871;
  assign T1827 = T1828 & RouterBuffer_5_io_deq_valid;
  assign T1828 = T1829 & T877;
  assign T1829 = T941 & T1830;
  assign T1830 = VCRouterStateManagement_5_io_currentState == 3'h4;
  assign T1831 = T1832 & T1824;
  assign T1832 = T1833 ^ 1'h1;
  assign T1833 = T943 | T951;
  assign readyToXmit_6_4 = T1834;
  assign T1834 = T1848 ? T1844 : T1835;
  assign T1835 = T1840 ? T1836 : 1'h0;
  assign T1836 = T1837 & RouterBuffer_6_io_deq_valid;
  assign T1837 = T1838 & T733;
  assign T1838 = T797 & T1839;
  assign T1839 = 3'h3 <= VCRouterStateManagement_6_io_currentState;
  assign T1840 = T806 & T1841;
  assign T1841 = T1842[3'h4:3'h4];
  assign T1842 = 1'h1 << T1843;
  assign T1843 = R727;
  assign T1844 = T1845 & RouterBuffer_6_io_deq_valid;
  assign T1845 = T1846 & T733;
  assign T1846 = T797 & T1847;
  assign T1847 = VCRouterStateManagement_6_io_currentState == 3'h4;
  assign T1848 = T1849 & T1841;
  assign T1849 = T1850 ^ 1'h1;
  assign T1850 = T799 | T807;
  assign readyToXmit_7_4 = T1851;
  assign T1851 = T1865 ? T1861 : T1852;
  assign T1852 = T1857 ? T1853 : 1'h0;
  assign T1853 = T1854 & RouterBuffer_7_io_deq_valid;
  assign T1854 = T1855 & T589;
  assign T1855 = T653 & T1856;
  assign T1856 = 3'h3 <= VCRouterStateManagement_7_io_currentState;
  assign T1857 = T662 & T1858;
  assign T1858 = T1859[3'h4:3'h4];
  assign T1859 = 1'h1 << T1860;
  assign T1860 = R583;
  assign T1861 = T1862 & RouterBuffer_7_io_deq_valid;
  assign T1862 = T1863 & T589;
  assign T1863 = T653 & T1864;
  assign T1864 = VCRouterStateManagement_7_io_currentState == 3'h4;
  assign T1865 = T1866 & T1858;
  assign T1866 = T1867 ^ 1'h1;
  assign T1867 = T655 | T663;
  assign T1868 = {readyToXmit_9_4, readyToXmit_8_4};
  assign readyToXmit_8_4 = T1869;
  assign T1869 = T1883 ? T1879 : T1870;
  assign T1870 = T1875 ? T1871 : 1'h0;
  assign T1871 = T1872 & RouterBuffer_8_io_deq_valid;
  assign T1872 = T1873 & T445;
  assign T1873 = T509 & T1874;
  assign T1874 = 3'h3 <= VCRouterStateManagement_8_io_currentState;
  assign T1875 = T518 & T1876;
  assign T1876 = T1877[3'h4:3'h4];
  assign T1877 = 1'h1 << T1878;
  assign T1878 = R439;
  assign T1879 = T1880 & RouterBuffer_8_io_deq_valid;
  assign T1880 = T1881 & T445;
  assign T1881 = T509 & T1882;
  assign T1882 = VCRouterStateManagement_8_io_currentState == 3'h4;
  assign T1883 = T1884 & T1876;
  assign T1884 = T1885 ^ 1'h1;
  assign T1885 = T511 | T519;
  assign readyToXmit_9_4 = T1886;
  assign T1886 = T1900 ? T1896 : T1887;
  assign T1887 = T1892 ? T1888 : 1'h0;
  assign T1888 = T1889 & RouterBuffer_9_io_deq_valid;
  assign T1889 = T1890 & T301;
  assign T1890 = T365 & T1891;
  assign T1891 = 3'h3 <= VCRouterStateManagement_9_io_currentState;
  assign T1892 = T374 & T1893;
  assign T1893 = T1894[3'h4:3'h4];
  assign T1894 = 1'h1 << T1895;
  assign T1895 = R295;
  assign T1896 = T1897 & RouterBuffer_9_io_deq_valid;
  assign T1897 = T1898 & T301;
  assign T1898 = T365 & T1899;
  assign T1899 = VCRouterStateManagement_9_io_currentState == 3'h4;
  assign T1900 = T1901 & T1893;
  assign T1901 = T1902 ^ 1'h1;
  assign T1902 = T367 | T375;
  assign T1903 = T1904 ? CreditCon_7_io_outCredit : CreditCon_6_io_outCredit;
  assign T1904 = T234;
  assign T1905 = T1906 != 10'h0;
  assign T1906 = T1907;
  assign T1907 = {T1937, T1908};
  assign T1908 = {T1926, T1909};
  assign T1909 = {readyToXmit_2_3, T1910};
  assign T1910 = {readyToXmit_1_3, readyToXmit_0_3};
  assign readyToXmit_0_3 = T1911;
  assign T1911 = T1915 ? T1738 : T1912;
  assign T1912 = T1913 ? T1730 : 1'h0;
  assign T1913 = T1670 & T1914;
  assign T1914 = T1736[2'h3:2'h3];
  assign T1915 = T1743 & T1914;
  assign readyToXmit_1_3 = T1916;
  assign T1916 = T1920 ? T1755 : T1917;
  assign T1917 = T1918 ? T1747 : 1'h0;
  assign T1918 = T1526 & T1919;
  assign T1919 = T1753[2'h3:2'h3];
  assign T1920 = T1760 & T1919;
  assign readyToXmit_2_3 = T1921;
  assign T1921 = T1925 ? T1772 : T1922;
  assign T1922 = T1923 ? T1764 : 1'h0;
  assign T1923 = T1382 & T1924;
  assign T1924 = T1770[2'h3:2'h3];
  assign T1925 = T1777 & T1924;
  assign T1926 = {readyToXmit_4_3, readyToXmit_3_3};
  assign readyToXmit_3_3 = T1927;
  assign T1927 = T1931 ? T1790 : T1928;
  assign T1928 = T1929 ? T1782 : 1'h0;
  assign T1929 = T1238 & T1930;
  assign T1930 = T1788[2'h3:2'h3];
  assign T1931 = T1795 & T1930;
  assign readyToXmit_4_3 = T1932;
  assign T1932 = T1936 ? T1807 : T1933;
  assign T1933 = T1934 ? T1799 : 1'h0;
  assign T1934 = T1094 & T1935;
  assign T1935 = T1805[2'h3:2'h3];
  assign T1936 = T1812 & T1935;
  assign T1937 = {T1955, T1938};
  assign T1938 = {readyToXmit_7_3, T1939};
  assign T1939 = {readyToXmit_6_3, readyToXmit_5_3};
  assign readyToXmit_5_3 = T1940;
  assign T1940 = T1944 ? T1827 : T1941;
  assign T1941 = T1942 ? T1819 : 1'h0;
  assign T1942 = T950 & T1943;
  assign T1943 = T1825[2'h3:2'h3];
  assign T1944 = T1832 & T1943;
  assign readyToXmit_6_3 = T1945;
  assign T1945 = T1949 ? T1844 : T1946;
  assign T1946 = T1947 ? T1836 : 1'h0;
  assign T1947 = T806 & T1948;
  assign T1948 = T1842[2'h3:2'h3];
  assign T1949 = T1849 & T1948;
  assign readyToXmit_7_3 = T1950;
  assign T1950 = T1954 ? T1861 : T1951;
  assign T1951 = T1952 ? T1853 : 1'h0;
  assign T1952 = T662 & T1953;
  assign T1953 = T1859[2'h3:2'h3];
  assign T1954 = T1866 & T1953;
  assign T1955 = {readyToXmit_9_3, readyToXmit_8_3};
  assign readyToXmit_8_3 = T1956;
  assign T1956 = T1960 ? T1879 : T1957;
  assign T1957 = T1958 ? T1871 : 1'h0;
  assign T1958 = T518 & T1959;
  assign T1959 = T1877[2'h3:2'h3];
  assign T1960 = T1884 & T1959;
  assign readyToXmit_9_3 = T1961;
  assign T1961 = T1965 ? T1896 : T1962;
  assign T1962 = T1963 ? T1888 : 1'h0;
  assign T1963 = T374 & T1964;
  assign T1964 = T1894[2'h3:2'h3];
  assign T1965 = T1901 & T1964;
  assign T1966 = T1967 ? CreditCon_5_io_outCredit : CreditCon_4_io_outCredit;
  assign T1967 = T246;
  assign T1968 = T1969 != 10'h0;
  assign T1969 = T1970;
  assign T1970 = {T2000, T1971};
  assign T1971 = {T1989, T1972};
  assign T1972 = {readyToXmit_2_2, T1973};
  assign T1973 = {readyToXmit_1_2, readyToXmit_0_2};
  assign readyToXmit_0_2 = T1974;
  assign T1974 = T1978 ? T1738 : T1975;
  assign T1975 = T1976 ? T1730 : 1'h0;
  assign T1976 = T1670 & T1977;
  assign T1977 = T1736[2'h2:2'h2];
  assign T1978 = T1743 & T1977;
  assign readyToXmit_1_2 = T1979;
  assign T1979 = T1983 ? T1755 : T1980;
  assign T1980 = T1981 ? T1747 : 1'h0;
  assign T1981 = T1526 & T1982;
  assign T1982 = T1753[2'h2:2'h2];
  assign T1983 = T1760 & T1982;
  assign readyToXmit_2_2 = T1984;
  assign T1984 = T1988 ? T1772 : T1985;
  assign T1985 = T1986 ? T1764 : 1'h0;
  assign T1986 = T1382 & T1987;
  assign T1987 = T1770[2'h2:2'h2];
  assign T1988 = T1777 & T1987;
  assign T1989 = {readyToXmit_4_2, readyToXmit_3_2};
  assign readyToXmit_3_2 = T1990;
  assign T1990 = T1994 ? T1790 : T1991;
  assign T1991 = T1992 ? T1782 : 1'h0;
  assign T1992 = T1238 & T1993;
  assign T1993 = T1788[2'h2:2'h2];
  assign T1994 = T1795 & T1993;
  assign readyToXmit_4_2 = T1995;
  assign T1995 = T1999 ? T1807 : T1996;
  assign T1996 = T1997 ? T1799 : 1'h0;
  assign T1997 = T1094 & T1998;
  assign T1998 = T1805[2'h2:2'h2];
  assign T1999 = T1812 & T1998;
  assign T2000 = {T2018, T2001};
  assign T2001 = {readyToXmit_7_2, T2002};
  assign T2002 = {readyToXmit_6_2, readyToXmit_5_2};
  assign readyToXmit_5_2 = T2003;
  assign T2003 = T2007 ? T1827 : T2004;
  assign T2004 = T2005 ? T1819 : 1'h0;
  assign T2005 = T950 & T2006;
  assign T2006 = T1825[2'h2:2'h2];
  assign T2007 = T1832 & T2006;
  assign readyToXmit_6_2 = T2008;
  assign T2008 = T2012 ? T1844 : T2009;
  assign T2009 = T2010 ? T1836 : 1'h0;
  assign T2010 = T806 & T2011;
  assign T2011 = T1842[2'h2:2'h2];
  assign T2012 = T1849 & T2011;
  assign readyToXmit_7_2 = T2013;
  assign T2013 = T2017 ? T1861 : T2014;
  assign T2014 = T2015 ? T1853 : 1'h0;
  assign T2015 = T662 & T2016;
  assign T2016 = T1859[2'h2:2'h2];
  assign T2017 = T1866 & T2016;
  assign T2018 = {readyToXmit_9_2, readyToXmit_8_2};
  assign readyToXmit_8_2 = T2019;
  assign T2019 = T2023 ? T1879 : T2020;
  assign T2020 = T2021 ? T1871 : 1'h0;
  assign T2021 = T518 & T2022;
  assign T2022 = T1877[2'h2:2'h2];
  assign T2023 = T1884 & T2022;
  assign readyToXmit_9_2 = T2024;
  assign T2024 = T2028 ? T1896 : T2025;
  assign T2025 = T2026 ? T1888 : 1'h0;
  assign T2026 = T374 & T2027;
  assign T2027 = T1894[2'h2:2'h2];
  assign T2028 = T1901 & T2027;
  assign T2029 = T2030 ? CreditCon_3_io_outCredit : CreditCon_2_io_outCredit;
  assign T2030 = T258;
  assign T2031 = T2032 != 10'h0;
  assign T2032 = T2033;
  assign T2033 = {T2063, T2034};
  assign T2034 = {T2052, T2035};
  assign T2035 = {readyToXmit_2_1, T2036};
  assign T2036 = {readyToXmit_1_1, readyToXmit_0_1};
  assign readyToXmit_0_1 = T2037;
  assign T2037 = T2041 ? T1738 : T2038;
  assign T2038 = T2039 ? T1730 : 1'h0;
  assign T2039 = T1670 & T2040;
  assign T2040 = T1736[1'h1:1'h1];
  assign T2041 = T1743 & T2040;
  assign readyToXmit_1_1 = T2042;
  assign T2042 = T2046 ? T1755 : T2043;
  assign T2043 = T2044 ? T1747 : 1'h0;
  assign T2044 = T1526 & T2045;
  assign T2045 = T1753[1'h1:1'h1];
  assign T2046 = T1760 & T2045;
  assign readyToXmit_2_1 = T2047;
  assign T2047 = T2051 ? T1772 : T2048;
  assign T2048 = T2049 ? T1764 : 1'h0;
  assign T2049 = T1382 & T2050;
  assign T2050 = T1770[1'h1:1'h1];
  assign T2051 = T1777 & T2050;
  assign T2052 = {readyToXmit_4_1, readyToXmit_3_1};
  assign readyToXmit_3_1 = T2053;
  assign T2053 = T2057 ? T1790 : T2054;
  assign T2054 = T2055 ? T1782 : 1'h0;
  assign T2055 = T1238 & T2056;
  assign T2056 = T1788[1'h1:1'h1];
  assign T2057 = T1795 & T2056;
  assign readyToXmit_4_1 = T2058;
  assign T2058 = T2062 ? T1807 : T2059;
  assign T2059 = T2060 ? T1799 : 1'h0;
  assign T2060 = T1094 & T2061;
  assign T2061 = T1805[1'h1:1'h1];
  assign T2062 = T1812 & T2061;
  assign T2063 = {T2081, T2064};
  assign T2064 = {readyToXmit_7_1, T2065};
  assign T2065 = {readyToXmit_6_1, readyToXmit_5_1};
  assign readyToXmit_5_1 = T2066;
  assign T2066 = T2070 ? T1827 : T2067;
  assign T2067 = T2068 ? T1819 : 1'h0;
  assign T2068 = T950 & T2069;
  assign T2069 = T1825[1'h1:1'h1];
  assign T2070 = T1832 & T2069;
  assign readyToXmit_6_1 = T2071;
  assign T2071 = T2075 ? T1844 : T2072;
  assign T2072 = T2073 ? T1836 : 1'h0;
  assign T2073 = T806 & T2074;
  assign T2074 = T1842[1'h1:1'h1];
  assign T2075 = T1849 & T2074;
  assign readyToXmit_7_1 = T2076;
  assign T2076 = T2080 ? T1861 : T2077;
  assign T2077 = T2078 ? T1853 : 1'h0;
  assign T2078 = T662 & T2079;
  assign T2079 = T1859[1'h1:1'h1];
  assign T2080 = T1866 & T2079;
  assign T2081 = {readyToXmit_9_1, readyToXmit_8_1};
  assign readyToXmit_8_1 = T2082;
  assign T2082 = T2086 ? T1879 : T2083;
  assign T2083 = T2084 ? T1871 : 1'h0;
  assign T2084 = T518 & T2085;
  assign T2085 = T1877[1'h1:1'h1];
  assign T2086 = T1884 & T2085;
  assign readyToXmit_9_1 = T2087;
  assign T2087 = T2091 ? T1896 : T2088;
  assign T2088 = T2089 ? T1888 : 1'h0;
  assign T2089 = T374 & T2090;
  assign T2090 = T1894[1'h1:1'h1];
  assign T2091 = T1901 & T2090;
  assign T2092 = T2093 ? CreditCon_1_io_outCredit : CreditCon_io_outCredit;
  assign T2093 = T270;
  assign T2094 = T2095 != 10'h0;
  assign T2095 = T2096;
  assign T2096 = {T2126, T2097};
  assign T2097 = {T2115, T2098};
  assign T2098 = {readyToXmit_2_0, T2099};
  assign T2099 = {readyToXmit_1_0, readyToXmit_0_0};
  assign readyToXmit_0_0 = T2100;
  assign T2100 = T2104 ? T1738 : T2101;
  assign T2101 = T2102 ? T1730 : 1'h0;
  assign T2102 = T1670 & T2103;
  assign T2103 = T1736[1'h0:1'h0];
  assign T2104 = T1743 & T2103;
  assign readyToXmit_1_0 = T2105;
  assign T2105 = T2109 ? T1755 : T2106;
  assign T2106 = T2107 ? T1747 : 1'h0;
  assign T2107 = T1526 & T2108;
  assign T2108 = T1753[1'h0:1'h0];
  assign T2109 = T1760 & T2108;
  assign readyToXmit_2_0 = T2110;
  assign T2110 = T2114 ? T1772 : T2111;
  assign T2111 = T2112 ? T1764 : 1'h0;
  assign T2112 = T1382 & T2113;
  assign T2113 = T1770[1'h0:1'h0];
  assign T2114 = T1777 & T2113;
  assign T2115 = {readyToXmit_4_0, readyToXmit_3_0};
  assign readyToXmit_3_0 = T2116;
  assign T2116 = T2120 ? T1790 : T2117;
  assign T2117 = T2118 ? T1782 : 1'h0;
  assign T2118 = T1238 & T2119;
  assign T2119 = T1788[1'h0:1'h0];
  assign T2120 = T1795 & T2119;
  assign readyToXmit_4_0 = T2121;
  assign T2121 = T2125 ? T1807 : T2122;
  assign T2122 = T2123 ? T1799 : 1'h0;
  assign T2123 = T1094 & T2124;
  assign T2124 = T1805[1'h0:1'h0];
  assign T2125 = T1812 & T2124;
  assign T2126 = {T2144, T2127};
  assign T2127 = {readyToXmit_7_0, T2128};
  assign T2128 = {readyToXmit_6_0, readyToXmit_5_0};
  assign readyToXmit_5_0 = T2129;
  assign T2129 = T2133 ? T1827 : T2130;
  assign T2130 = T2131 ? T1819 : 1'h0;
  assign T2131 = T950 & T2132;
  assign T2132 = T1825[1'h0:1'h0];
  assign T2133 = T1832 & T2132;
  assign readyToXmit_6_0 = T2134;
  assign T2134 = T2138 ? T1844 : T2135;
  assign T2135 = T2136 ? T1836 : 1'h0;
  assign T2136 = T806 & T2137;
  assign T2137 = T1842[1'h0:1'h0];
  assign T2138 = T1849 & T2137;
  assign readyToXmit_7_0 = T2139;
  assign T2139 = T2143 ? T1861 : T2140;
  assign T2140 = T2141 ? T1853 : 1'h0;
  assign T2141 = T662 & T2142;
  assign T2142 = T1859[1'h0:1'h0];
  assign T2143 = T1866 & T2142;
  assign T2144 = {readyToXmit_9_0, readyToXmit_8_0};
  assign readyToXmit_8_0 = T2145;
  assign T2145 = T2149 ? T1879 : T2146;
  assign T2146 = T2147 ? T1871 : 1'h0;
  assign T2147 = T518 & T2148;
  assign T2148 = T1877[1'h0:1'h0];
  assign T2149 = T1884 & T2148;
  assign readyToXmit_9_0 = T2150;
  assign T2150 = T2154 ? T1896 : T2151;
  assign T2151 = T2152 ? T1888 : 1'h0;
  assign T2152 = T374 & T2153;
  assign T2153 = T1894[1'h0:1'h0];
  assign T2154 = T1901 & T2153;
  assign T2155 = RouterBuffer_io_deq_valid & T2156;
  assign T2156 = 3'h2 <= VCRouterStateManagement_io_currentState;
  assign T2157 = RouterBuffer_1_io_deq_valid & T2158;
  assign T2158 = 3'h2 <= VCRouterStateManagement_1_io_currentState;
  assign T2159 = RouterBuffer_2_io_deq_valid & T2160;
  assign T2160 = 3'h2 <= VCRouterStateManagement_2_io_currentState;
  assign T2161 = RouterBuffer_3_io_deq_valid & T2162;
  assign T2162 = 3'h2 <= VCRouterStateManagement_3_io_currentState;
  assign T2163 = RouterBuffer_4_io_deq_valid & T2164;
  assign T2164 = 3'h2 <= VCRouterStateManagement_4_io_currentState;
  assign T2165 = RouterBuffer_5_io_deq_valid & T2166;
  assign T2166 = 3'h2 <= VCRouterStateManagement_5_io_currentState;
  assign T2167 = RouterBuffer_6_io_deq_valid & T2168;
  assign T2168 = 3'h2 <= VCRouterStateManagement_6_io_currentState;
  assign T2169 = RouterBuffer_7_io_deq_valid & T2170;
  assign T2170 = 3'h2 <= VCRouterStateManagement_7_io_currentState;
  assign T2171 = RouterBuffer_8_io_deq_valid & T2172;
  assign T2172 = 3'h2 <= VCRouterStateManagement_8_io_currentState;
  assign T2173 = RouterBuffer_9_io_deq_valid & T2174;
  assign T2174 = 3'h2 <= VCRouterStateManagement_9_io_currentState;
  assign T2175 = validVCs_0_0[1'h0:1'h0];
  assign T2177 = T2179 & T2178;
  assign T2178 = VCRouterOutputStateManagement_io_currentState == 2'h2;
  assign T2179 = flitsAreTail_0 & CreditCon_io_outCredit;
  assign T2180 = validVCs_0_0[1'h1:1'h1];
  assign T2182 = T2184 & T2183;
  assign T2183 = VCRouterOutputStateManagement_io_currentState == 2'h2;
  assign T2184 = flitsAreTail_0 & CreditCon_1_io_outCredit;
  assign T2185 = validVCs_0_1[1'h0:1'h0];
  assign T2187 = T2189 & T2188;
  assign T2188 = VCRouterOutputStateManagement_1_io_currentState == 2'h2;
  assign T2189 = flitsAreTail_0 & CreditCon_2_io_outCredit;
  assign T2190 = validVCs_0_1[1'h1:1'h1];
  assign T2192 = T2194 & T2193;
  assign T2193 = VCRouterOutputStateManagement_1_io_currentState == 2'h2;
  assign T2194 = flitsAreTail_0 & CreditCon_3_io_outCredit;
  assign T2195 = validVCs_0_2[1'h0:1'h0];
  assign T2197 = T2199 & T2198;
  assign T2198 = VCRouterOutputStateManagement_2_io_currentState == 2'h2;
  assign T2199 = flitsAreTail_0 & CreditCon_4_io_outCredit;
  assign T2200 = validVCs_0_2[1'h1:1'h1];
  assign T2202 = T2204 & T2203;
  assign T2203 = VCRouterOutputStateManagement_2_io_currentState == 2'h2;
  assign T2204 = flitsAreTail_0 & CreditCon_5_io_outCredit;
  assign T2205 = validVCs_0_3[1'h0:1'h0];
  assign T2207 = T2209 & T2208;
  assign T2208 = VCRouterOutputStateManagement_3_io_currentState == 2'h2;
  assign T2209 = flitsAreTail_0 & CreditCon_6_io_outCredit;
  assign T2210 = validVCs_0_3[1'h1:1'h1];
  assign T2212 = T2214 & T2213;
  assign T2213 = VCRouterOutputStateManagement_3_io_currentState == 2'h2;
  assign T2214 = flitsAreTail_0 & CreditCon_7_io_outCredit;
  assign T2215 = validVCs_0_4[1'h0:1'h0];
  assign T2217 = T2219 & T2218;
  assign T2218 = VCRouterOutputStateManagement_4_io_currentState == 2'h2;
  assign T2219 = flitsAreTail_0 & CreditCon_8_io_outCredit;
  assign T2220 = validVCs_0_4[1'h1:1'h1];
  assign T2222 = T2224 & T2223;
  assign T2223 = VCRouterOutputStateManagement_4_io_currentState == 2'h2;
  assign T2224 = flitsAreTail_0 & CreditCon_9_io_outCredit;
  assign T2225 = validVCs_1_0[1'h0:1'h0];
  assign T2227 = T2229 & T2228;
  assign T2228 = VCRouterOutputStateManagement_io_currentState == 2'h2;
  assign T2229 = flitsAreTail_1 & CreditCon_io_outCredit;
  assign T2230 = validVCs_1_0[1'h1:1'h1];
  assign T2232 = T2234 & T2233;
  assign T2233 = VCRouterOutputStateManagement_io_currentState == 2'h2;
  assign T2234 = flitsAreTail_1 & CreditCon_1_io_outCredit;
  assign T2235 = validVCs_1_1[1'h0:1'h0];
  assign T2237 = T2239 & T2238;
  assign T2238 = VCRouterOutputStateManagement_1_io_currentState == 2'h2;
  assign T2239 = flitsAreTail_1 & CreditCon_2_io_outCredit;
  assign T2240 = validVCs_1_1[1'h1:1'h1];
  assign T2242 = T2244 & T2243;
  assign T2243 = VCRouterOutputStateManagement_1_io_currentState == 2'h2;
  assign T2244 = flitsAreTail_1 & CreditCon_3_io_outCredit;
  assign T2245 = validVCs_1_2[1'h0:1'h0];
  assign T2247 = T2249 & T2248;
  assign T2248 = VCRouterOutputStateManagement_2_io_currentState == 2'h2;
  assign T2249 = flitsAreTail_1 & CreditCon_4_io_outCredit;
  assign T2250 = validVCs_1_2[1'h1:1'h1];
  assign T2252 = T2254 & T2253;
  assign T2253 = VCRouterOutputStateManagement_2_io_currentState == 2'h2;
  assign T2254 = flitsAreTail_1 & CreditCon_5_io_outCredit;
  assign T2255 = validVCs_1_3[1'h0:1'h0];
  assign T2257 = T2259 & T2258;
  assign T2258 = VCRouterOutputStateManagement_3_io_currentState == 2'h2;
  assign T2259 = flitsAreTail_1 & CreditCon_6_io_outCredit;
  assign T2260 = validVCs_1_3[1'h1:1'h1];
  assign T2262 = T2264 & T2263;
  assign T2263 = VCRouterOutputStateManagement_3_io_currentState == 2'h2;
  assign T2264 = flitsAreTail_1 & CreditCon_7_io_outCredit;
  assign T2265 = validVCs_1_4[1'h0:1'h0];
  assign T2267 = T2269 & T2268;
  assign T2268 = VCRouterOutputStateManagement_4_io_currentState == 2'h2;
  assign T2269 = flitsAreTail_1 & CreditCon_8_io_outCredit;
  assign T2270 = validVCs_1_4[1'h1:1'h1];
  assign T2272 = T2274 & T2273;
  assign T2273 = VCRouterOutputStateManagement_4_io_currentState == 2'h2;
  assign T2274 = flitsAreTail_1 & CreditCon_9_io_outCredit;
  assign T2275 = validVCs_2_0[1'h0:1'h0];
  assign T2277 = T2279 & T2278;
  assign T2278 = VCRouterOutputStateManagement_io_currentState == 2'h2;
  assign T2279 = flitsAreTail_2 & CreditCon_io_outCredit;
  assign T2280 = validVCs_2_0[1'h1:1'h1];
  assign T2282 = T2284 & T2283;
  assign T2283 = VCRouterOutputStateManagement_io_currentState == 2'h2;
  assign T2284 = flitsAreTail_2 & CreditCon_1_io_outCredit;
  assign T2285 = validVCs_2_1[1'h0:1'h0];
  assign T2287 = T2289 & T2288;
  assign T2288 = VCRouterOutputStateManagement_1_io_currentState == 2'h2;
  assign T2289 = flitsAreTail_2 & CreditCon_2_io_outCredit;
  assign T2290 = validVCs_2_1[1'h1:1'h1];
  assign T2292 = T2294 & T2293;
  assign T2293 = VCRouterOutputStateManagement_1_io_currentState == 2'h2;
  assign T2294 = flitsAreTail_2 & CreditCon_3_io_outCredit;
  assign T2295 = validVCs_2_2[1'h0:1'h0];
  assign T2297 = T2299 & T2298;
  assign T2298 = VCRouterOutputStateManagement_2_io_currentState == 2'h2;
  assign T2299 = flitsAreTail_2 & CreditCon_4_io_outCredit;
  assign T2300 = validVCs_2_2[1'h1:1'h1];
  assign T2302 = T2304 & T2303;
  assign T2303 = VCRouterOutputStateManagement_2_io_currentState == 2'h2;
  assign T2304 = flitsAreTail_2 & CreditCon_5_io_outCredit;
  assign T2305 = validVCs_2_3[1'h0:1'h0];
  assign T2307 = T2309 & T2308;
  assign T2308 = VCRouterOutputStateManagement_3_io_currentState == 2'h2;
  assign T2309 = flitsAreTail_2 & CreditCon_6_io_outCredit;
  assign T2310 = validVCs_2_3[1'h1:1'h1];
  assign T2312 = T2314 & T2313;
  assign T2313 = VCRouterOutputStateManagement_3_io_currentState == 2'h2;
  assign T2314 = flitsAreTail_2 & CreditCon_7_io_outCredit;
  assign T2315 = validVCs_2_4[1'h0:1'h0];
  assign T2317 = T2319 & T2318;
  assign T2318 = VCRouterOutputStateManagement_4_io_currentState == 2'h2;
  assign T2319 = flitsAreTail_2 & CreditCon_8_io_outCredit;
  assign T2320 = validVCs_2_4[1'h1:1'h1];
  assign T2322 = T2324 & T2323;
  assign T2323 = VCRouterOutputStateManagement_4_io_currentState == 2'h2;
  assign T2324 = flitsAreTail_2 & CreditCon_9_io_outCredit;
  assign T2325 = validVCs_3_0[1'h0:1'h0];
  assign T2327 = T2329 & T2328;
  assign T2328 = VCRouterOutputStateManagement_io_currentState == 2'h2;
  assign T2329 = flitsAreTail_3 & CreditCon_io_outCredit;
  assign T2330 = validVCs_3_0[1'h1:1'h1];
  assign T2332 = T2334 & T2333;
  assign T2333 = VCRouterOutputStateManagement_io_currentState == 2'h2;
  assign T2334 = flitsAreTail_3 & CreditCon_1_io_outCredit;
  assign T2335 = validVCs_3_1[1'h0:1'h0];
  assign T2337 = T2339 & T2338;
  assign T2338 = VCRouterOutputStateManagement_1_io_currentState == 2'h2;
  assign T2339 = flitsAreTail_3 & CreditCon_2_io_outCredit;
  assign T2340 = validVCs_3_1[1'h1:1'h1];
  assign T2342 = T2344 & T2343;
  assign T2343 = VCRouterOutputStateManagement_1_io_currentState == 2'h2;
  assign T2344 = flitsAreTail_3 & CreditCon_3_io_outCredit;
  assign T2345 = validVCs_3_2[1'h0:1'h0];
  assign T2347 = T2349 & T2348;
  assign T2348 = VCRouterOutputStateManagement_2_io_currentState == 2'h2;
  assign T2349 = flitsAreTail_3 & CreditCon_4_io_outCredit;
  assign T2350 = validVCs_3_2[1'h1:1'h1];
  assign T2352 = T2354 & T2353;
  assign T2353 = VCRouterOutputStateManagement_2_io_currentState == 2'h2;
  assign T2354 = flitsAreTail_3 & CreditCon_5_io_outCredit;
  assign T2355 = validVCs_3_3[1'h0:1'h0];
  assign T2357 = T2359 & T2358;
  assign T2358 = VCRouterOutputStateManagement_3_io_currentState == 2'h2;
  assign T2359 = flitsAreTail_3 & CreditCon_6_io_outCredit;
  assign T2360 = validVCs_3_3[1'h1:1'h1];
  assign T2362 = T2364 & T2363;
  assign T2363 = VCRouterOutputStateManagement_3_io_currentState == 2'h2;
  assign T2364 = flitsAreTail_3 & CreditCon_7_io_outCredit;
  assign T2365 = validVCs_3_4[1'h0:1'h0];
  assign T2367 = T2369 & T2368;
  assign T2368 = VCRouterOutputStateManagement_4_io_currentState == 2'h2;
  assign T2369 = flitsAreTail_3 & CreditCon_8_io_outCredit;
  assign T2370 = validVCs_3_4[1'h1:1'h1];
  assign T2372 = T2374 & T2373;
  assign T2373 = VCRouterOutputStateManagement_4_io_currentState == 2'h2;
  assign T2374 = flitsAreTail_3 & CreditCon_9_io_outCredit;
  assign T2375 = validVCs_4_0[1'h0:1'h0];
  assign T2377 = T2379 & T2378;
  assign T2378 = VCRouterOutputStateManagement_io_currentState == 2'h2;
  assign T2379 = flitsAreTail_4 & CreditCon_io_outCredit;
  assign T2380 = validVCs_4_0[1'h1:1'h1];
  assign T2382 = T2384 & T2383;
  assign T2383 = VCRouterOutputStateManagement_io_currentState == 2'h2;
  assign T2384 = flitsAreTail_4 & CreditCon_1_io_outCredit;
  assign T2385 = validVCs_4_1[1'h0:1'h0];
  assign T2387 = T2389 & T2388;
  assign T2388 = VCRouterOutputStateManagement_1_io_currentState == 2'h2;
  assign T2389 = flitsAreTail_4 & CreditCon_2_io_outCredit;
  assign T2390 = validVCs_4_1[1'h1:1'h1];
  assign T2392 = T2394 & T2393;
  assign T2393 = VCRouterOutputStateManagement_1_io_currentState == 2'h2;
  assign T2394 = flitsAreTail_4 & CreditCon_3_io_outCredit;
  assign T2395 = validVCs_4_2[1'h0:1'h0];
  assign T2397 = T2399 & T2398;
  assign T2398 = VCRouterOutputStateManagement_2_io_currentState == 2'h2;
  assign T2399 = flitsAreTail_4 & CreditCon_4_io_outCredit;
  assign T2400 = validVCs_4_2[1'h1:1'h1];
  assign T2402 = T2404 & T2403;
  assign T2403 = VCRouterOutputStateManagement_2_io_currentState == 2'h2;
  assign T2404 = flitsAreTail_4 & CreditCon_5_io_outCredit;
  assign T2405 = validVCs_4_3[1'h0:1'h0];
  assign T2407 = T2409 & T2408;
  assign T2408 = VCRouterOutputStateManagement_3_io_currentState == 2'h2;
  assign T2409 = flitsAreTail_4 & CreditCon_6_io_outCredit;
  assign T2410 = validVCs_4_3[1'h1:1'h1];
  assign T2412 = T2414 & T2413;
  assign T2413 = VCRouterOutputStateManagement_3_io_currentState == 2'h2;
  assign T2414 = flitsAreTail_4 & CreditCon_7_io_outCredit;
  assign T2415 = validVCs_4_4[1'h0:1'h0];
  assign T2417 = T2419 & T2418;
  assign T2418 = VCRouterOutputStateManagement_4_io_currentState == 2'h2;
  assign T2419 = flitsAreTail_4 & CreditCon_8_io_outCredit;
  assign T2420 = validVCs_4_4[1'h1:1'h1];
  assign T2422 = T2424 & T2423;
  assign T2423 = VCRouterOutputStateManagement_4_io_currentState == 2'h2;
  assign T2424 = flitsAreTail_4 & CreditCon_9_io_outCredit;
  assign T2425 = validVCs_5_0[1'h0:1'h0];
  assign T2427 = T2429 & T2428;
  assign T2428 = VCRouterOutputStateManagement_io_currentState == 2'h2;
  assign T2429 = flitsAreTail_5 & CreditCon_io_outCredit;
  assign T2430 = validVCs_5_0[1'h1:1'h1];
  assign T2432 = T2434 & T2433;
  assign T2433 = VCRouterOutputStateManagement_io_currentState == 2'h2;
  assign T2434 = flitsAreTail_5 & CreditCon_1_io_outCredit;
  assign T2435 = validVCs_5_1[1'h0:1'h0];
  assign T2437 = T2439 & T2438;
  assign T2438 = VCRouterOutputStateManagement_1_io_currentState == 2'h2;
  assign T2439 = flitsAreTail_5 & CreditCon_2_io_outCredit;
  assign T2440 = validVCs_5_1[1'h1:1'h1];
  assign T2442 = T2444 & T2443;
  assign T2443 = VCRouterOutputStateManagement_1_io_currentState == 2'h2;
  assign T2444 = flitsAreTail_5 & CreditCon_3_io_outCredit;
  assign T2445 = validVCs_5_2[1'h0:1'h0];
  assign T2447 = T2449 & T2448;
  assign T2448 = VCRouterOutputStateManagement_2_io_currentState == 2'h2;
  assign T2449 = flitsAreTail_5 & CreditCon_4_io_outCredit;
  assign T2450 = validVCs_5_2[1'h1:1'h1];
  assign T2452 = T2454 & T2453;
  assign T2453 = VCRouterOutputStateManagement_2_io_currentState == 2'h2;
  assign T2454 = flitsAreTail_5 & CreditCon_5_io_outCredit;
  assign T2455 = validVCs_5_3[1'h0:1'h0];
  assign T2457 = T2459 & T2458;
  assign T2458 = VCRouterOutputStateManagement_3_io_currentState == 2'h2;
  assign T2459 = flitsAreTail_5 & CreditCon_6_io_outCredit;
  assign T2460 = validVCs_5_3[1'h1:1'h1];
  assign T2462 = T2464 & T2463;
  assign T2463 = VCRouterOutputStateManagement_3_io_currentState == 2'h2;
  assign T2464 = flitsAreTail_5 & CreditCon_7_io_outCredit;
  assign T2465 = validVCs_5_4[1'h0:1'h0];
  assign T2467 = T2469 & T2468;
  assign T2468 = VCRouterOutputStateManagement_4_io_currentState == 2'h2;
  assign T2469 = flitsAreTail_5 & CreditCon_8_io_outCredit;
  assign T2470 = validVCs_5_4[1'h1:1'h1];
  assign T2472 = T2474 & T2473;
  assign T2473 = VCRouterOutputStateManagement_4_io_currentState == 2'h2;
  assign T2474 = flitsAreTail_5 & CreditCon_9_io_outCredit;
  assign T2475 = validVCs_6_0[1'h0:1'h0];
  assign T2477 = T2479 & T2478;
  assign T2478 = VCRouterOutputStateManagement_io_currentState == 2'h2;
  assign T2479 = flitsAreTail_6 & CreditCon_io_outCredit;
  assign T2480 = validVCs_6_0[1'h1:1'h1];
  assign T2482 = T2484 & T2483;
  assign T2483 = VCRouterOutputStateManagement_io_currentState == 2'h2;
  assign T2484 = flitsAreTail_6 & CreditCon_1_io_outCredit;
  assign T2485 = validVCs_6_1[1'h0:1'h0];
  assign T2487 = T2489 & T2488;
  assign T2488 = VCRouterOutputStateManagement_1_io_currentState == 2'h2;
  assign T2489 = flitsAreTail_6 & CreditCon_2_io_outCredit;
  assign T2490 = validVCs_6_1[1'h1:1'h1];
  assign T2492 = T2494 & T2493;
  assign T2493 = VCRouterOutputStateManagement_1_io_currentState == 2'h2;
  assign T2494 = flitsAreTail_6 & CreditCon_3_io_outCredit;
  assign T2495 = validVCs_6_2[1'h0:1'h0];
  assign T2497 = T2499 & T2498;
  assign T2498 = VCRouterOutputStateManagement_2_io_currentState == 2'h2;
  assign T2499 = flitsAreTail_6 & CreditCon_4_io_outCredit;
  assign T2500 = validVCs_6_2[1'h1:1'h1];
  assign T2502 = T2504 & T2503;
  assign T2503 = VCRouterOutputStateManagement_2_io_currentState == 2'h2;
  assign T2504 = flitsAreTail_6 & CreditCon_5_io_outCredit;
  assign T2505 = validVCs_6_3[1'h0:1'h0];
  assign T2507 = T2509 & T2508;
  assign T2508 = VCRouterOutputStateManagement_3_io_currentState == 2'h2;
  assign T2509 = flitsAreTail_6 & CreditCon_6_io_outCredit;
  assign T2510 = validVCs_6_3[1'h1:1'h1];
  assign T2512 = T2514 & T2513;
  assign T2513 = VCRouterOutputStateManagement_3_io_currentState == 2'h2;
  assign T2514 = flitsAreTail_6 & CreditCon_7_io_outCredit;
  assign T2515 = validVCs_6_4[1'h0:1'h0];
  assign T2517 = T2519 & T2518;
  assign T2518 = VCRouterOutputStateManagement_4_io_currentState == 2'h2;
  assign T2519 = flitsAreTail_6 & CreditCon_8_io_outCredit;
  assign T2520 = validVCs_6_4[1'h1:1'h1];
  assign T2522 = T2524 & T2523;
  assign T2523 = VCRouterOutputStateManagement_4_io_currentState == 2'h2;
  assign T2524 = flitsAreTail_6 & CreditCon_9_io_outCredit;
  assign T2525 = validVCs_7_0[1'h0:1'h0];
  assign T2527 = T2529 & T2528;
  assign T2528 = VCRouterOutputStateManagement_io_currentState == 2'h2;
  assign T2529 = flitsAreTail_7 & CreditCon_io_outCredit;
  assign T2530 = validVCs_7_0[1'h1:1'h1];
  assign T2532 = T2534 & T2533;
  assign T2533 = VCRouterOutputStateManagement_io_currentState == 2'h2;
  assign T2534 = flitsAreTail_7 & CreditCon_1_io_outCredit;
  assign T2535 = validVCs_7_1[1'h0:1'h0];
  assign T2537 = T2539 & T2538;
  assign T2538 = VCRouterOutputStateManagement_1_io_currentState == 2'h2;
  assign T2539 = flitsAreTail_7 & CreditCon_2_io_outCredit;
  assign T2540 = validVCs_7_1[1'h1:1'h1];
  assign T2542 = T2544 & T2543;
  assign T2543 = VCRouterOutputStateManagement_1_io_currentState == 2'h2;
  assign T2544 = flitsAreTail_7 & CreditCon_3_io_outCredit;
  assign T2545 = validVCs_7_2[1'h0:1'h0];
  assign T2547 = T2549 & T2548;
  assign T2548 = VCRouterOutputStateManagement_2_io_currentState == 2'h2;
  assign T2549 = flitsAreTail_7 & CreditCon_4_io_outCredit;
  assign T2550 = validVCs_7_2[1'h1:1'h1];
  assign T2552 = T2554 & T2553;
  assign T2553 = VCRouterOutputStateManagement_2_io_currentState == 2'h2;
  assign T2554 = flitsAreTail_7 & CreditCon_5_io_outCredit;
  assign T2555 = validVCs_7_3[1'h0:1'h0];
  assign T2557 = T2559 & T2558;
  assign T2558 = VCRouterOutputStateManagement_3_io_currentState == 2'h2;
  assign T2559 = flitsAreTail_7 & CreditCon_6_io_outCredit;
  assign T2560 = validVCs_7_3[1'h1:1'h1];
  assign T2562 = T2564 & T2563;
  assign T2563 = VCRouterOutputStateManagement_3_io_currentState == 2'h2;
  assign T2564 = flitsAreTail_7 & CreditCon_7_io_outCredit;
  assign T2565 = validVCs_7_4[1'h0:1'h0];
  assign T2567 = T2569 & T2568;
  assign T2568 = VCRouterOutputStateManagement_4_io_currentState == 2'h2;
  assign T2569 = flitsAreTail_7 & CreditCon_8_io_outCredit;
  assign T2570 = validVCs_7_4[1'h1:1'h1];
  assign T2572 = T2574 & T2573;
  assign T2573 = VCRouterOutputStateManagement_4_io_currentState == 2'h2;
  assign T2574 = flitsAreTail_7 & CreditCon_9_io_outCredit;
  assign T2575 = validVCs_8_0[1'h0:1'h0];
  assign T2577 = T2579 & T2578;
  assign T2578 = VCRouterOutputStateManagement_io_currentState == 2'h2;
  assign T2579 = flitsAreTail_8 & CreditCon_io_outCredit;
  assign T2580 = validVCs_8_0[1'h1:1'h1];
  assign T2582 = T2584 & T2583;
  assign T2583 = VCRouterOutputStateManagement_io_currentState == 2'h2;
  assign T2584 = flitsAreTail_8 & CreditCon_1_io_outCredit;
  assign T2585 = validVCs_8_1[1'h0:1'h0];
  assign T2587 = T2589 & T2588;
  assign T2588 = VCRouterOutputStateManagement_1_io_currentState == 2'h2;
  assign T2589 = flitsAreTail_8 & CreditCon_2_io_outCredit;
  assign T2590 = validVCs_8_1[1'h1:1'h1];
  assign T2592 = T2594 & T2593;
  assign T2593 = VCRouterOutputStateManagement_1_io_currentState == 2'h2;
  assign T2594 = flitsAreTail_8 & CreditCon_3_io_outCredit;
  assign T2595 = validVCs_8_2[1'h0:1'h0];
  assign T2597 = T2599 & T2598;
  assign T2598 = VCRouterOutputStateManagement_2_io_currentState == 2'h2;
  assign T2599 = flitsAreTail_8 & CreditCon_4_io_outCredit;
  assign T2600 = validVCs_8_2[1'h1:1'h1];
  assign T2602 = T2604 & T2603;
  assign T2603 = VCRouterOutputStateManagement_2_io_currentState == 2'h2;
  assign T2604 = flitsAreTail_8 & CreditCon_5_io_outCredit;
  assign T2605 = validVCs_8_3[1'h0:1'h0];
  assign T2607 = T2609 & T2608;
  assign T2608 = VCRouterOutputStateManagement_3_io_currentState == 2'h2;
  assign T2609 = flitsAreTail_8 & CreditCon_6_io_outCredit;
  assign T2610 = validVCs_8_3[1'h1:1'h1];
  assign T2612 = T2614 & T2613;
  assign T2613 = VCRouterOutputStateManagement_3_io_currentState == 2'h2;
  assign T2614 = flitsAreTail_8 & CreditCon_7_io_outCredit;
  assign T2615 = validVCs_8_4[1'h0:1'h0];
  assign T2617 = T2619 & T2618;
  assign T2618 = VCRouterOutputStateManagement_4_io_currentState == 2'h2;
  assign T2619 = flitsAreTail_8 & CreditCon_8_io_outCredit;
  assign T2620 = validVCs_8_4[1'h1:1'h1];
  assign T2622 = T2624 & T2623;
  assign T2623 = VCRouterOutputStateManagement_4_io_currentState == 2'h2;
  assign T2624 = flitsAreTail_8 & CreditCon_9_io_outCredit;
  assign T2625 = validVCs_9_0[1'h0:1'h0];
  assign T2627 = T2629 & T2628;
  assign T2628 = VCRouterOutputStateManagement_io_currentState == 2'h2;
  assign T2629 = flitsAreTail_9 & CreditCon_io_outCredit;
  assign T2630 = validVCs_9_0[1'h1:1'h1];
  assign T2632 = T2634 & T2633;
  assign T2633 = VCRouterOutputStateManagement_io_currentState == 2'h2;
  assign T2634 = flitsAreTail_9 & CreditCon_1_io_outCredit;
  assign T2635 = validVCs_9_1[1'h0:1'h0];
  assign T2637 = T2639 & T2638;
  assign T2638 = VCRouterOutputStateManagement_1_io_currentState == 2'h2;
  assign T2639 = flitsAreTail_9 & CreditCon_2_io_outCredit;
  assign T2640 = validVCs_9_1[1'h1:1'h1];
  assign T2642 = T2644 & T2643;
  assign T2643 = VCRouterOutputStateManagement_1_io_currentState == 2'h2;
  assign T2644 = flitsAreTail_9 & CreditCon_3_io_outCredit;
  assign T2645 = validVCs_9_2[1'h0:1'h0];
  assign T2647 = T2649 & T2648;
  assign T2648 = VCRouterOutputStateManagement_2_io_currentState == 2'h2;
  assign T2649 = flitsAreTail_9 & CreditCon_4_io_outCredit;
  assign T2650 = validVCs_9_2[1'h1:1'h1];
  assign T2652 = T2654 & T2653;
  assign T2653 = VCRouterOutputStateManagement_2_io_currentState == 2'h2;
  assign T2654 = flitsAreTail_9 & CreditCon_5_io_outCredit;
  assign T2655 = validVCs_9_3[1'h0:1'h0];
  assign T2657 = T2659 & T2658;
  assign T2658 = VCRouterOutputStateManagement_3_io_currentState == 2'h2;
  assign T2659 = flitsAreTail_9 & CreditCon_6_io_outCredit;
  assign T2660 = validVCs_9_3[1'h1:1'h1];
  assign T2662 = T2664 & T2663;
  assign T2663 = VCRouterOutputStateManagement_3_io_currentState == 2'h2;
  assign T2664 = flitsAreTail_9 & CreditCon_7_io_outCredit;
  assign T2665 = validVCs_9_4[1'h0:1'h0];
  assign T2667 = T2669 & T2668;
  assign T2668 = VCRouterOutputStateManagement_4_io_currentState == 2'h2;
  assign T2669 = flitsAreTail_9 & CreditCon_8_io_outCredit;
  assign T2670 = validVCs_9_4[1'h1:1'h1];
  assign T2672 = T2674 & T2673;
  assign T2673 = VCRouterOutputStateManagement_4_io_currentState == 2'h2;
  assign T2674 = flitsAreTail_9 & CreditCon_9_io_outCredit;
  assign T3182 = reset ? 3'h0 : T2676;
  assign T2676 = T1670 ? T2677 : R2675;
  assign T2677 = T2678[2'h2:1'h0];
  assign T2678 = RouterBuffer_io_deq_bits_x[5'h1f:1'h1];
  assign T2679 = T2681 & T2680;
  assign T2680 = 3'h3 <= VCRouterStateManagement_io_currentState;
  assign T2681 = T2682;
  assign T2682 = R2683[1'h0:1'h0];
  assign T3183 = reset ? 8'h0 : T2684;
  assign T2684 = 1'h1 << CMeshDOR_io_result;
  assign T2685 = T2687 & T2686;
  assign T2686 = VCRouterStateManagement_io_currentState == 3'h4;
  assign T2687 = R2688;
  assign T3184 = reset ? 1'h1 : T1692;
  assign T3185 = reset ? 3'h0 : T2690;
  assign T2690 = T1526 ? T2691 : R2689;
  assign T2691 = T2692[2'h2:1'h0];
  assign T2692 = RouterBuffer_1_io_deq_bits_x[5'h1f:1'h1];
  assign T2693 = T2695 & T2694;
  assign T2694 = 3'h3 <= VCRouterStateManagement_1_io_currentState;
  assign T2695 = T2696;
  assign T2696 = R2697[1'h0:1'h0];
  assign T3186 = reset ? 8'h0 : T2698;
  assign T2698 = 1'h1 << CMeshDOR_1_io_result;
  assign T2699 = T2701 & T2700;
  assign T2700 = VCRouterStateManagement_1_io_currentState == 3'h4;
  assign T2701 = R2702;
  assign T3187 = reset ? 1'h1 : T1548;
  assign T3188 = reset ? 3'h0 : T2704;
  assign T2704 = T1382 ? T2705 : R2703;
  assign T2705 = T2706[2'h2:1'h0];
  assign T2706 = RouterBuffer_2_io_deq_bits_x[5'h1f:1'h1];
  assign T2707 = T2709 & T2708;
  assign T2708 = 3'h3 <= VCRouterStateManagement_2_io_currentState;
  assign T2709 = T2710;
  assign T2710 = R2711[1'h0:1'h0];
  assign T3189 = reset ? 8'h0 : T2712;
  assign T2712 = 1'h1 << CMeshDOR_2_io_result;
  assign T2713 = T2715 & T2714;
  assign T2714 = VCRouterStateManagement_2_io_currentState == 3'h4;
  assign T2715 = R2716;
  assign T3190 = reset ? 1'h1 : T1404;
  assign T3191 = reset ? 3'h0 : T2718;
  assign T2718 = T1238 ? T2719 : R2717;
  assign T2719 = T2720[2'h2:1'h0];
  assign T2720 = RouterBuffer_3_io_deq_bits_x[5'h1f:1'h1];
  assign T2721 = T2723 & T2722;
  assign T2722 = 3'h3 <= VCRouterStateManagement_3_io_currentState;
  assign T2723 = T2724;
  assign T2724 = R2725[1'h0:1'h0];
  assign T3192 = reset ? 8'h0 : T2726;
  assign T2726 = 1'h1 << CMeshDOR_3_io_result;
  assign T2727 = T2729 & T2728;
  assign T2728 = VCRouterStateManagement_3_io_currentState == 3'h4;
  assign T2729 = R2730;
  assign T3193 = reset ? 1'h1 : T1260;
  assign T3194 = reset ? 3'h0 : T2732;
  assign T2732 = T1094 ? T2733 : R2731;
  assign T2733 = T2734[2'h2:1'h0];
  assign T2734 = RouterBuffer_4_io_deq_bits_x[5'h1f:1'h1];
  assign T2735 = T2737 & T2736;
  assign T2736 = 3'h3 <= VCRouterStateManagement_4_io_currentState;
  assign T2737 = T2738;
  assign T2738 = R2739[1'h0:1'h0];
  assign T3195 = reset ? 8'h0 : T2740;
  assign T2740 = 1'h1 << CMeshDOR_4_io_result;
  assign T2741 = T2743 & T2742;
  assign T2742 = VCRouterStateManagement_4_io_currentState == 3'h4;
  assign T2743 = R2744;
  assign T3196 = reset ? 1'h1 : T1116;
  assign T3197 = reset ? 3'h0 : T2746;
  assign T2746 = T950 ? T2747 : R2745;
  assign T2747 = T2748[2'h2:1'h0];
  assign T2748 = RouterBuffer_5_io_deq_bits_x[5'h1f:1'h1];
  assign T2749 = T2751 & T2750;
  assign T2750 = 3'h3 <= VCRouterStateManagement_5_io_currentState;
  assign T2751 = T2752;
  assign T2752 = R2753[1'h0:1'h0];
  assign T3198 = reset ? 8'h0 : T2754;
  assign T2754 = 1'h1 << CMeshDOR_5_io_result;
  assign T2755 = T2757 & T2756;
  assign T2756 = VCRouterStateManagement_5_io_currentState == 3'h4;
  assign T2757 = R2758;
  assign T3199 = reset ? 1'h1 : T972;
  assign T3200 = reset ? 3'h0 : T2760;
  assign T2760 = T806 ? T2761 : R2759;
  assign T2761 = T2762[2'h2:1'h0];
  assign T2762 = RouterBuffer_6_io_deq_bits_x[5'h1f:1'h1];
  assign T2763 = T2765 & T2764;
  assign T2764 = 3'h3 <= VCRouterStateManagement_6_io_currentState;
  assign T2765 = T2766;
  assign T2766 = R2767[1'h0:1'h0];
  assign T3201 = reset ? 8'h0 : T2768;
  assign T2768 = 1'h1 << CMeshDOR_6_io_result;
  assign T2769 = T2771 & T2770;
  assign T2770 = VCRouterStateManagement_6_io_currentState == 3'h4;
  assign T2771 = R2772;
  assign T3202 = reset ? 1'h1 : T828;
  assign T3203 = reset ? 3'h0 : T2774;
  assign T2774 = T662 ? T2775 : R2773;
  assign T2775 = T2776[2'h2:1'h0];
  assign T2776 = RouterBuffer_7_io_deq_bits_x[5'h1f:1'h1];
  assign T2777 = T2779 & T2778;
  assign T2778 = 3'h3 <= VCRouterStateManagement_7_io_currentState;
  assign T2779 = T2780;
  assign T2780 = R2781[1'h0:1'h0];
  assign T3204 = reset ? 8'h0 : T2782;
  assign T2782 = 1'h1 << CMeshDOR_7_io_result;
  assign T2783 = T2785 & T2784;
  assign T2784 = VCRouterStateManagement_7_io_currentState == 3'h4;
  assign T2785 = R2786;
  assign T3205 = reset ? 1'h1 : T684;
  assign T3206 = reset ? 3'h0 : T2788;
  assign T2788 = T518 ? T2789 : R2787;
  assign T2789 = T2790[2'h2:1'h0];
  assign T2790 = RouterBuffer_8_io_deq_bits_x[5'h1f:1'h1];
  assign T2791 = T2793 & T2792;
  assign T2792 = 3'h3 <= VCRouterStateManagement_8_io_currentState;
  assign T2793 = T2794;
  assign T2794 = R2795[1'h0:1'h0];
  assign T3207 = reset ? 8'h0 : T2796;
  assign T2796 = 1'h1 << CMeshDOR_8_io_result;
  assign T2797 = T2799 & T2798;
  assign T2798 = VCRouterStateManagement_8_io_currentState == 3'h4;
  assign T2799 = R2800;
  assign T3208 = reset ? 1'h1 : T540;
  assign T3209 = reset ? 3'h0 : T2802;
  assign T2802 = T374 ? T2803 : R2801;
  assign T2803 = T2804[2'h2:1'h0];
  assign T2804 = RouterBuffer_9_io_deq_bits_x[5'h1f:1'h1];
  assign T2805 = T2807 & T2806;
  assign T2806 = 3'h3 <= VCRouterStateManagement_9_io_currentState;
  assign T2807 = T2808;
  assign T2808 = R2809[1'h0:1'h0];
  assign T3210 = reset ? 8'h0 : T2810;
  assign T2810 = 1'h1 << CMeshDOR_9_io_result;
  assign T2811 = T2813 & T2812;
  assign T2812 = VCRouterStateManagement_9_io_currentState == 3'h4;
  assign T2813 = R2814;
  assign T3211 = reset ? 1'h1 : T396;
  assign T2815 = T2817 & T2816;
  assign T2816 = 3'h3 <= VCRouterStateManagement_io_currentState;
  assign T2817 = T2818;
  assign T2818 = R2683[1'h1:1'h1];
  assign T2819 = T2821 & T2820;
  assign T2820 = VCRouterStateManagement_io_currentState == 3'h4;
  assign T2821 = R2688;
  assign T2822 = T2824 & T2823;
  assign T2823 = 3'h3 <= VCRouterStateManagement_1_io_currentState;
  assign T2824 = T2825;
  assign T2825 = R2697[1'h1:1'h1];
  assign T2826 = T2828 & T2827;
  assign T2827 = VCRouterStateManagement_1_io_currentState == 3'h4;
  assign T2828 = R2702;
  assign T2829 = T2831 & T2830;
  assign T2830 = 3'h3 <= VCRouterStateManagement_2_io_currentState;
  assign T2831 = T2832;
  assign T2832 = R2711[1'h1:1'h1];
  assign T2833 = T2835 & T2834;
  assign T2834 = VCRouterStateManagement_2_io_currentState == 3'h4;
  assign T2835 = R2716;
  assign T2836 = T2838 & T2837;
  assign T2837 = 3'h3 <= VCRouterStateManagement_3_io_currentState;
  assign T2838 = T2839;
  assign T2839 = R2725[1'h1:1'h1];
  assign T2840 = T2842 & T2841;
  assign T2841 = VCRouterStateManagement_3_io_currentState == 3'h4;
  assign T2842 = R2730;
  assign T2843 = T2845 & T2844;
  assign T2844 = 3'h3 <= VCRouterStateManagement_4_io_currentState;
  assign T2845 = T2846;
  assign T2846 = R2739[1'h1:1'h1];
  assign T2847 = T2849 & T2848;
  assign T2848 = VCRouterStateManagement_4_io_currentState == 3'h4;
  assign T2849 = R2744;
  assign T2850 = T2852 & T2851;
  assign T2851 = 3'h3 <= VCRouterStateManagement_5_io_currentState;
  assign T2852 = T2853;
  assign T2853 = R2753[1'h1:1'h1];
  assign T2854 = T2856 & T2855;
  assign T2855 = VCRouterStateManagement_5_io_currentState == 3'h4;
  assign T2856 = R2758;
  assign T2857 = T2859 & T2858;
  assign T2858 = 3'h3 <= VCRouterStateManagement_6_io_currentState;
  assign T2859 = T2860;
  assign T2860 = R2767[1'h1:1'h1];
  assign T2861 = T2863 & T2862;
  assign T2862 = VCRouterStateManagement_6_io_currentState == 3'h4;
  assign T2863 = R2772;
  assign T2864 = T2866 & T2865;
  assign T2865 = 3'h3 <= VCRouterStateManagement_7_io_currentState;
  assign T2866 = T2867;
  assign T2867 = R2781[1'h1:1'h1];
  assign T2868 = T2870 & T2869;
  assign T2869 = VCRouterStateManagement_7_io_currentState == 3'h4;
  assign T2870 = R2786;
  assign T2871 = T2873 & T2872;
  assign T2872 = 3'h3 <= VCRouterStateManagement_8_io_currentState;
  assign T2873 = T2874;
  assign T2874 = R2795[1'h1:1'h1];
  assign T2875 = T2877 & T2876;
  assign T2876 = VCRouterStateManagement_8_io_currentState == 3'h4;
  assign T2877 = R2800;
  assign T2878 = T2880 & T2879;
  assign T2879 = 3'h3 <= VCRouterStateManagement_9_io_currentState;
  assign T2880 = T2881;
  assign T2881 = R2809[1'h1:1'h1];
  assign T2882 = T2884 & T2883;
  assign T2883 = VCRouterStateManagement_9_io_currentState == 3'h4;
  assign T2884 = R2814;
  assign T2885 = T2887 & T2886;
  assign T2886 = 3'h3 <= VCRouterStateManagement_io_currentState;
  assign T2887 = T2888;
  assign T2888 = R2683[2'h2:2'h2];
  assign T2889 = T2891 & T2890;
  assign T2890 = VCRouterStateManagement_io_currentState == 3'h4;
  assign T2891 = R2688;
  assign T2892 = T2894 & T2893;
  assign T2893 = 3'h3 <= VCRouterStateManagement_1_io_currentState;
  assign T2894 = T2895;
  assign T2895 = R2697[2'h2:2'h2];
  assign T2896 = T2898 & T2897;
  assign T2897 = VCRouterStateManagement_1_io_currentState == 3'h4;
  assign T2898 = R2702;
  assign T2899 = T2901 & T2900;
  assign T2900 = 3'h3 <= VCRouterStateManagement_2_io_currentState;
  assign T2901 = T2902;
  assign T2902 = R2711[2'h2:2'h2];
  assign T2903 = T2905 & T2904;
  assign T2904 = VCRouterStateManagement_2_io_currentState == 3'h4;
  assign T2905 = R2716;
  assign T2906 = T2908 & T2907;
  assign T2907 = 3'h3 <= VCRouterStateManagement_3_io_currentState;
  assign T2908 = T2909;
  assign T2909 = R2725[2'h2:2'h2];
  assign T2910 = T2912 & T2911;
  assign T2911 = VCRouterStateManagement_3_io_currentState == 3'h4;
  assign T2912 = R2730;
  assign T2913 = T2915 & T2914;
  assign T2914 = 3'h3 <= VCRouterStateManagement_4_io_currentState;
  assign T2915 = T2916;
  assign T2916 = R2739[2'h2:2'h2];
  assign T2917 = T2919 & T2918;
  assign T2918 = VCRouterStateManagement_4_io_currentState == 3'h4;
  assign T2919 = R2744;
  assign T2920 = T2922 & T2921;
  assign T2921 = 3'h3 <= VCRouterStateManagement_5_io_currentState;
  assign T2922 = T2923;
  assign T2923 = R2753[2'h2:2'h2];
  assign T2924 = T2926 & T2925;
  assign T2925 = VCRouterStateManagement_5_io_currentState == 3'h4;
  assign T2926 = R2758;
  assign T2927 = T2929 & T2928;
  assign T2928 = 3'h3 <= VCRouterStateManagement_6_io_currentState;
  assign T2929 = T2930;
  assign T2930 = R2767[2'h2:2'h2];
  assign T2931 = T2933 & T2932;
  assign T2932 = VCRouterStateManagement_6_io_currentState == 3'h4;
  assign T2933 = R2772;
  assign T2934 = T2936 & T2935;
  assign T2935 = 3'h3 <= VCRouterStateManagement_7_io_currentState;
  assign T2936 = T2937;
  assign T2937 = R2781[2'h2:2'h2];
  assign T2938 = T2940 & T2939;
  assign T2939 = VCRouterStateManagement_7_io_currentState == 3'h4;
  assign T2940 = R2786;
  assign T2941 = T2943 & T2942;
  assign T2942 = 3'h3 <= VCRouterStateManagement_8_io_currentState;
  assign T2943 = T2944;
  assign T2944 = R2795[2'h2:2'h2];
  assign T2945 = T2947 & T2946;
  assign T2946 = VCRouterStateManagement_8_io_currentState == 3'h4;
  assign T2947 = R2800;
  assign T2948 = T2950 & T2949;
  assign T2949 = 3'h3 <= VCRouterStateManagement_9_io_currentState;
  assign T2950 = T2951;
  assign T2951 = R2809[2'h2:2'h2];
  assign T2952 = T2954 & T2953;
  assign T2953 = VCRouterStateManagement_9_io_currentState == 3'h4;
  assign T2954 = R2814;
  assign T2955 = T2957 & T2956;
  assign T2956 = 3'h3 <= VCRouterStateManagement_io_currentState;
  assign T2957 = T2958;
  assign T2958 = R2683[2'h3:2'h3];
  assign T2959 = T2961 & T2960;
  assign T2960 = VCRouterStateManagement_io_currentState == 3'h4;
  assign T2961 = R2688;
  assign T2962 = T2964 & T2963;
  assign T2963 = 3'h3 <= VCRouterStateManagement_1_io_currentState;
  assign T2964 = T2965;
  assign T2965 = R2697[2'h3:2'h3];
  assign T2966 = T2968 & T2967;
  assign T2967 = VCRouterStateManagement_1_io_currentState == 3'h4;
  assign T2968 = R2702;
  assign T2969 = T2971 & T2970;
  assign T2970 = 3'h3 <= VCRouterStateManagement_2_io_currentState;
  assign T2971 = T2972;
  assign T2972 = R2711[2'h3:2'h3];
  assign T2973 = T2975 & T2974;
  assign T2974 = VCRouterStateManagement_2_io_currentState == 3'h4;
  assign T2975 = R2716;
  assign T2976 = T2978 & T2977;
  assign T2977 = 3'h3 <= VCRouterStateManagement_3_io_currentState;
  assign T2978 = T2979;
  assign T2979 = R2725[2'h3:2'h3];
  assign T2980 = T2982 & T2981;
  assign T2981 = VCRouterStateManagement_3_io_currentState == 3'h4;
  assign T2982 = R2730;
  assign T2983 = T2985 & T2984;
  assign T2984 = 3'h3 <= VCRouterStateManagement_4_io_currentState;
  assign T2985 = T2986;
  assign T2986 = R2739[2'h3:2'h3];
  assign T2987 = T2989 & T2988;
  assign T2988 = VCRouterStateManagement_4_io_currentState == 3'h4;
  assign T2989 = R2744;
  assign T2990 = T2992 & T2991;
  assign T2991 = 3'h3 <= VCRouterStateManagement_5_io_currentState;
  assign T2992 = T2993;
  assign T2993 = R2753[2'h3:2'h3];
  assign T2994 = T2996 & T2995;
  assign T2995 = VCRouterStateManagement_5_io_currentState == 3'h4;
  assign T2996 = R2758;
  assign T2997 = T2999 & T2998;
  assign T2998 = 3'h3 <= VCRouterStateManagement_6_io_currentState;
  assign T2999 = T3000;
  assign T3000 = R2767[2'h3:2'h3];
  assign T3001 = T3003 & T3002;
  assign T3002 = VCRouterStateManagement_6_io_currentState == 3'h4;
  assign T3003 = R2772;
  assign T3004 = T3006 & T3005;
  assign T3005 = 3'h3 <= VCRouterStateManagement_7_io_currentState;
  assign T3006 = T3007;
  assign T3007 = R2781[2'h3:2'h3];
  assign T3008 = T3010 & T3009;
  assign T3009 = VCRouterStateManagement_7_io_currentState == 3'h4;
  assign T3010 = R2786;
  assign T3011 = T3013 & T3012;
  assign T3012 = 3'h3 <= VCRouterStateManagement_8_io_currentState;
  assign T3013 = T3014;
  assign T3014 = R2795[2'h3:2'h3];
  assign T3015 = T3017 & T3016;
  assign T3016 = VCRouterStateManagement_8_io_currentState == 3'h4;
  assign T3017 = R2800;
  assign T3018 = T3020 & T3019;
  assign T3019 = 3'h3 <= VCRouterStateManagement_9_io_currentState;
  assign T3020 = T3021;
  assign T3021 = R2809[2'h3:2'h3];
  assign T3022 = T3024 & T3023;
  assign T3023 = VCRouterStateManagement_9_io_currentState == 3'h4;
  assign T3024 = R2814;
  assign T3025 = T3027 & T3026;
  assign T3026 = 3'h3 <= VCRouterStateManagement_io_currentState;
  assign T3027 = T3028;
  assign T3028 = R2683[3'h4:3'h4];
  assign T3029 = T3031 & T3030;
  assign T3030 = VCRouterStateManagement_io_currentState == 3'h4;
  assign T3031 = R2688;
  assign T3032 = T3034 & T3033;
  assign T3033 = 3'h3 <= VCRouterStateManagement_1_io_currentState;
  assign T3034 = T3035;
  assign T3035 = R2697[3'h4:3'h4];
  assign T3036 = T3038 & T3037;
  assign T3037 = VCRouterStateManagement_1_io_currentState == 3'h4;
  assign T3038 = R2702;
  assign T3039 = T3041 & T3040;
  assign T3040 = 3'h3 <= VCRouterStateManagement_2_io_currentState;
  assign T3041 = T3042;
  assign T3042 = R2711[3'h4:3'h4];
  assign T3043 = T3045 & T3044;
  assign T3044 = VCRouterStateManagement_2_io_currentState == 3'h4;
  assign T3045 = R2716;
  assign T3046 = T3048 & T3047;
  assign T3047 = 3'h3 <= VCRouterStateManagement_3_io_currentState;
  assign T3048 = T3049;
  assign T3049 = R2725[3'h4:3'h4];
  assign T3050 = T3052 & T3051;
  assign T3051 = VCRouterStateManagement_3_io_currentState == 3'h4;
  assign T3052 = R2730;
  assign T3053 = T3055 & T3054;
  assign T3054 = 3'h3 <= VCRouterStateManagement_4_io_currentState;
  assign T3055 = T3056;
  assign T3056 = R2739[3'h4:3'h4];
  assign T3057 = T3059 & T3058;
  assign T3058 = VCRouterStateManagement_4_io_currentState == 3'h4;
  assign T3059 = R2744;
  assign T3060 = T3062 & T3061;
  assign T3061 = 3'h3 <= VCRouterStateManagement_5_io_currentState;
  assign T3062 = T3063;
  assign T3063 = R2753[3'h4:3'h4];
  assign T3064 = T3066 & T3065;
  assign T3065 = VCRouterStateManagement_5_io_currentState == 3'h4;
  assign T3066 = R2758;
  assign T3067 = T3069 & T3068;
  assign T3068 = 3'h3 <= VCRouterStateManagement_6_io_currentState;
  assign T3069 = T3070;
  assign T3070 = R2767[3'h4:3'h4];
  assign T3071 = T3073 & T3072;
  assign T3072 = VCRouterStateManagement_6_io_currentState == 3'h4;
  assign T3073 = R2772;
  assign T3074 = T3076 & T3075;
  assign T3075 = 3'h3 <= VCRouterStateManagement_7_io_currentState;
  assign T3076 = T3077;
  assign T3077 = R2781[3'h4:3'h4];
  assign T3078 = T3080 & T3079;
  assign T3079 = VCRouterStateManagement_7_io_currentState == 3'h4;
  assign T3080 = R2786;
  assign T3081 = T3083 & T3082;
  assign T3082 = 3'h3 <= VCRouterStateManagement_8_io_currentState;
  assign T3083 = T3084;
  assign T3084 = R2795[3'h4:3'h4];
  assign T3085 = T3087 & T3086;
  assign T3086 = VCRouterStateManagement_8_io_currentState == 3'h4;
  assign T3087 = R2800;
  assign T3088 = T3090 & T3089;
  assign T3089 = 3'h3 <= VCRouterStateManagement_9_io_currentState;
  assign T3090 = T3091;
  assign T3091 = R2809[3'h4:3'h4];
  assign T3092 = T3094 & T3093;
  assign T3093 = VCRouterStateManagement_9_io_currentState == 3'h4;
  assign T3094 = R2814;
  assign io_counters_0_counterVal = T3212;
  assign T3212 = {31'h0, T3095};
  assign T3095 = T3096 == 1'h0;
  assign T3096 = T365 ^ 1'h1;
  assign io_outChannels_0_flitValid = R3097;
  assign io_outChannels_0_flit_x = R3098;
  assign T3099 = 55'h0;
  assign T3213 = reset ? T3099 : switch_io_outPorts_0_x;
  assign io_outChannels_1_flitValid = R3100;
  assign io_outChannels_1_flit_x = R3101;
  assign T3102 = 55'h0;
  assign T3214 = reset ? T3102 : switch_io_outPorts_1_x;
  assign io_outChannels_2_flitValid = R3103;
  assign io_outChannels_2_flit_x = R3104;
  assign T3105 = 55'h0;
  assign T3215 = reset ? T3105 : switch_io_outPorts_2_x;
  assign io_outChannels_3_flitValid = R3106;
  assign io_outChannels_3_flit_x = R3107;
  assign T3108 = 55'h0;
  assign T3216 = reset ? T3108 : switch_io_outPorts_3_x;
  assign io_outChannels_4_flitValid = R3109;
  assign io_outChannels_4_flit_x = R3110;
  assign T3111 = 55'h0;
  assign T3217 = reset ? T3111 : switch_io_outPorts_4_x;
  assign io_inChannels_0_credit_0_grant = CreditGen_io_outCredit_grant;
  assign io_inChannels_0_credit_1_grant = CreditGen_1_io_outCredit_grant;
  assign io_inChannels_1_credit_0_grant = CreditGen_2_io_outCredit_grant;
  assign io_inChannels_1_credit_1_grant = CreditGen_3_io_outCredit_grant;
  assign io_inChannels_2_credit_0_grant = CreditGen_4_io_outCredit_grant;
  assign io_inChannels_2_credit_1_grant = CreditGen_5_io_outCredit_grant;
  assign io_inChannels_3_credit_0_grant = CreditGen_6_io_outCredit_grant;
  assign io_inChannels_3_credit_1_grant = CreditGen_7_io_outCredit_grant;
  assign io_inChannels_4_credit_0_grant = CreditGen_8_io_outCredit_grant;
  assign io_inChannels_4_credit_1_grant = CreditGen_9_io_outCredit_grant;
  Switch switch(
       .io_inPorts_9_x( ReplaceVCPort_9_io_newFlit_x ),
       .io_inPorts_8_x( ReplaceVCPort_8_io_newFlit_x ),
       .io_inPorts_7_x( ReplaceVCPort_7_io_newFlit_x ),
       .io_inPorts_6_x( ReplaceVCPort_6_io_newFlit_x ),
       .io_inPorts_5_x( ReplaceVCPort_5_io_newFlit_x ),
       .io_inPorts_4_x( ReplaceVCPort_4_io_newFlit_x ),
       .io_inPorts_3_x( ReplaceVCPort_3_io_newFlit_x ),
       .io_inPorts_2_x( ReplaceVCPort_2_io_newFlit_x ),
       .io_inPorts_1_x( ReplaceVCPort_1_io_newFlit_x ),
       .io_inPorts_0_x( ReplaceVCPort_io_newFlit_x ),
       .io_outPorts_4_x( switch_io_outPorts_4_x ),
       .io_outPorts_3_x( switch_io_outPorts_3_x ),
       .io_outPorts_2_x( switch_io_outPorts_2_x ),
       .io_outPorts_1_x( switch_io_outPorts_1_x ),
       .io_outPorts_0_x( switch_io_outPorts_0_x ),
       .io_sel_4( swAllocator_io_chosens_4 ),
       .io_sel_3( swAllocator_io_chosens_3 ),
       .io_sel_2( swAllocator_io_chosens_2 ),
       .io_sel_1( swAllocator_io_chosens_1 ),
       .io_sel_0( swAllocator_io_chosens_0 )
  );
  SwitchAllocator_0 swAllocator(.clk(clk), .reset(reset),
       .io_requests_4_9_releaseLock( T3092 ),
       .io_requests_4_9_grant( swAllocator_io_requests_4_9_grant ),
       .io_requests_4_9_request( T3088 ),
       .io_requests_4_9_priorityLevel( R2801 ),
       .io_requests_4_8_releaseLock( T3085 ),
       .io_requests_4_8_grant( swAllocator_io_requests_4_8_grant ),
       .io_requests_4_8_request( T3081 ),
       .io_requests_4_8_priorityLevel( R2787 ),
       .io_requests_4_7_releaseLock( T3078 ),
       .io_requests_4_7_grant( swAllocator_io_requests_4_7_grant ),
       .io_requests_4_7_request( T3074 ),
       .io_requests_4_7_priorityLevel( R2773 ),
       .io_requests_4_6_releaseLock( T3071 ),
       .io_requests_4_6_grant( swAllocator_io_requests_4_6_grant ),
       .io_requests_4_6_request( T3067 ),
       .io_requests_4_6_priorityLevel( R2759 ),
       .io_requests_4_5_releaseLock( T3064 ),
       .io_requests_4_5_grant( swAllocator_io_requests_4_5_grant ),
       .io_requests_4_5_request( T3060 ),
       .io_requests_4_5_priorityLevel( R2745 ),
       .io_requests_4_4_releaseLock( T3057 ),
       .io_requests_4_4_grant( swAllocator_io_requests_4_4_grant ),
       .io_requests_4_4_request( T3053 ),
       .io_requests_4_4_priorityLevel( R2731 ),
       .io_requests_4_3_releaseLock( T3050 ),
       .io_requests_4_3_grant( swAllocator_io_requests_4_3_grant ),
       .io_requests_4_3_request( T3046 ),
       .io_requests_4_3_priorityLevel( R2717 ),
       .io_requests_4_2_releaseLock( T3043 ),
       .io_requests_4_2_grant( swAllocator_io_requests_4_2_grant ),
       .io_requests_4_2_request( T3039 ),
       .io_requests_4_2_priorityLevel( R2703 ),
       .io_requests_4_1_releaseLock( T3036 ),
       .io_requests_4_1_grant( swAllocator_io_requests_4_1_grant ),
       .io_requests_4_1_request( T3032 ),
       .io_requests_4_1_priorityLevel( R2689 ),
       .io_requests_4_0_releaseLock( T3029 ),
       .io_requests_4_0_grant( swAllocator_io_requests_4_0_grant ),
       .io_requests_4_0_request( T3025 ),
       .io_requests_4_0_priorityLevel( R2675 ),
       .io_requests_3_9_releaseLock( T3022 ),
       .io_requests_3_9_grant( swAllocator_io_requests_3_9_grant ),
       .io_requests_3_9_request( T3018 ),
       .io_requests_3_9_priorityLevel( R2801 ),
       .io_requests_3_8_releaseLock( T3015 ),
       .io_requests_3_8_grant( swAllocator_io_requests_3_8_grant ),
       .io_requests_3_8_request( T3011 ),
       .io_requests_3_8_priorityLevel( R2787 ),
       .io_requests_3_7_releaseLock( T3008 ),
       .io_requests_3_7_grant( swAllocator_io_requests_3_7_grant ),
       .io_requests_3_7_request( T3004 ),
       .io_requests_3_7_priorityLevel( R2773 ),
       .io_requests_3_6_releaseLock( T3001 ),
       .io_requests_3_6_grant( swAllocator_io_requests_3_6_grant ),
       .io_requests_3_6_request( T2997 ),
       .io_requests_3_6_priorityLevel( R2759 ),
       .io_requests_3_5_releaseLock( T2994 ),
       .io_requests_3_5_grant( swAllocator_io_requests_3_5_grant ),
       .io_requests_3_5_request( T2990 ),
       .io_requests_3_5_priorityLevel( R2745 ),
       .io_requests_3_4_releaseLock( T2987 ),
       .io_requests_3_4_grant( swAllocator_io_requests_3_4_grant ),
       .io_requests_3_4_request( T2983 ),
       .io_requests_3_4_priorityLevel( R2731 ),
       .io_requests_3_3_releaseLock( T2980 ),
       .io_requests_3_3_grant( swAllocator_io_requests_3_3_grant ),
       .io_requests_3_3_request( T2976 ),
       .io_requests_3_3_priorityLevel( R2717 ),
       .io_requests_3_2_releaseLock( T2973 ),
       .io_requests_3_2_grant( swAllocator_io_requests_3_2_grant ),
       .io_requests_3_2_request( T2969 ),
       .io_requests_3_2_priorityLevel( R2703 ),
       .io_requests_3_1_releaseLock( T2966 ),
       .io_requests_3_1_grant( swAllocator_io_requests_3_1_grant ),
       .io_requests_3_1_request( T2962 ),
       .io_requests_3_1_priorityLevel( R2689 ),
       .io_requests_3_0_releaseLock( T2959 ),
       .io_requests_3_0_grant( swAllocator_io_requests_3_0_grant ),
       .io_requests_3_0_request( T2955 ),
       .io_requests_3_0_priorityLevel( R2675 ),
       .io_requests_2_9_releaseLock( T2952 ),
       .io_requests_2_9_grant( swAllocator_io_requests_2_9_grant ),
       .io_requests_2_9_request( T2948 ),
       .io_requests_2_9_priorityLevel( R2801 ),
       .io_requests_2_8_releaseLock( T2945 ),
       .io_requests_2_8_grant( swAllocator_io_requests_2_8_grant ),
       .io_requests_2_8_request( T2941 ),
       .io_requests_2_8_priorityLevel( R2787 ),
       .io_requests_2_7_releaseLock( T2938 ),
       .io_requests_2_7_grant( swAllocator_io_requests_2_7_grant ),
       .io_requests_2_7_request( T2934 ),
       .io_requests_2_7_priorityLevel( R2773 ),
       .io_requests_2_6_releaseLock( T2931 ),
       .io_requests_2_6_grant( swAllocator_io_requests_2_6_grant ),
       .io_requests_2_6_request( T2927 ),
       .io_requests_2_6_priorityLevel( R2759 ),
       .io_requests_2_5_releaseLock( T2924 ),
       .io_requests_2_5_grant( swAllocator_io_requests_2_5_grant ),
       .io_requests_2_5_request( T2920 ),
       .io_requests_2_5_priorityLevel( R2745 ),
       .io_requests_2_4_releaseLock( T2917 ),
       .io_requests_2_4_grant( swAllocator_io_requests_2_4_grant ),
       .io_requests_2_4_request( T2913 ),
       .io_requests_2_4_priorityLevel( R2731 ),
       .io_requests_2_3_releaseLock( T2910 ),
       .io_requests_2_3_grant( swAllocator_io_requests_2_3_grant ),
       .io_requests_2_3_request( T2906 ),
       .io_requests_2_3_priorityLevel( R2717 ),
       .io_requests_2_2_releaseLock( T2903 ),
       .io_requests_2_2_grant( swAllocator_io_requests_2_2_grant ),
       .io_requests_2_2_request( T2899 ),
       .io_requests_2_2_priorityLevel( R2703 ),
       .io_requests_2_1_releaseLock( T2896 ),
       .io_requests_2_1_grant( swAllocator_io_requests_2_1_grant ),
       .io_requests_2_1_request( T2892 ),
       .io_requests_2_1_priorityLevel( R2689 ),
       .io_requests_2_0_releaseLock( T2889 ),
       .io_requests_2_0_grant( swAllocator_io_requests_2_0_grant ),
       .io_requests_2_0_request( T2885 ),
       .io_requests_2_0_priorityLevel( R2675 ),
       .io_requests_1_9_releaseLock( T2882 ),
       .io_requests_1_9_grant( swAllocator_io_requests_1_9_grant ),
       .io_requests_1_9_request( T2878 ),
       .io_requests_1_9_priorityLevel( R2801 ),
       .io_requests_1_8_releaseLock( T2875 ),
       .io_requests_1_8_grant( swAllocator_io_requests_1_8_grant ),
       .io_requests_1_8_request( T2871 ),
       .io_requests_1_8_priorityLevel( R2787 ),
       .io_requests_1_7_releaseLock( T2868 ),
       .io_requests_1_7_grant( swAllocator_io_requests_1_7_grant ),
       .io_requests_1_7_request( T2864 ),
       .io_requests_1_7_priorityLevel( R2773 ),
       .io_requests_1_6_releaseLock( T2861 ),
       .io_requests_1_6_grant( swAllocator_io_requests_1_6_grant ),
       .io_requests_1_6_request( T2857 ),
       .io_requests_1_6_priorityLevel( R2759 ),
       .io_requests_1_5_releaseLock( T2854 ),
       .io_requests_1_5_grant( swAllocator_io_requests_1_5_grant ),
       .io_requests_1_5_request( T2850 ),
       .io_requests_1_5_priorityLevel( R2745 ),
       .io_requests_1_4_releaseLock( T2847 ),
       .io_requests_1_4_grant( swAllocator_io_requests_1_4_grant ),
       .io_requests_1_4_request( T2843 ),
       .io_requests_1_4_priorityLevel( R2731 ),
       .io_requests_1_3_releaseLock( T2840 ),
       .io_requests_1_3_grant( swAllocator_io_requests_1_3_grant ),
       .io_requests_1_3_request( T2836 ),
       .io_requests_1_3_priorityLevel( R2717 ),
       .io_requests_1_2_releaseLock( T2833 ),
       .io_requests_1_2_grant( swAllocator_io_requests_1_2_grant ),
       .io_requests_1_2_request( T2829 ),
       .io_requests_1_2_priorityLevel( R2703 ),
       .io_requests_1_1_releaseLock( T2826 ),
       .io_requests_1_1_grant( swAllocator_io_requests_1_1_grant ),
       .io_requests_1_1_request( T2822 ),
       .io_requests_1_1_priorityLevel( R2689 ),
       .io_requests_1_0_releaseLock( T2819 ),
       .io_requests_1_0_grant( swAllocator_io_requests_1_0_grant ),
       .io_requests_1_0_request( T2815 ),
       .io_requests_1_0_priorityLevel( R2675 ),
       .io_requests_0_9_releaseLock( T2811 ),
       .io_requests_0_9_grant( swAllocator_io_requests_0_9_grant ),
       .io_requests_0_9_request( T2805 ),
       .io_requests_0_9_priorityLevel( R2801 ),
       .io_requests_0_8_releaseLock( T2797 ),
       .io_requests_0_8_grant( swAllocator_io_requests_0_8_grant ),
       .io_requests_0_8_request( T2791 ),
       .io_requests_0_8_priorityLevel( R2787 ),
       .io_requests_0_7_releaseLock( T2783 ),
       .io_requests_0_7_grant( swAllocator_io_requests_0_7_grant ),
       .io_requests_0_7_request( T2777 ),
       .io_requests_0_7_priorityLevel( R2773 ),
       .io_requests_0_6_releaseLock( T2769 ),
       .io_requests_0_6_grant( swAllocator_io_requests_0_6_grant ),
       .io_requests_0_6_request( T2763 ),
       .io_requests_0_6_priorityLevel( R2759 ),
       .io_requests_0_5_releaseLock( T2755 ),
       .io_requests_0_5_grant( swAllocator_io_requests_0_5_grant ),
       .io_requests_0_5_request( T2749 ),
       .io_requests_0_5_priorityLevel( R2745 ),
       .io_requests_0_4_releaseLock( T2741 ),
       .io_requests_0_4_grant( swAllocator_io_requests_0_4_grant ),
       .io_requests_0_4_request( T2735 ),
       .io_requests_0_4_priorityLevel( R2731 ),
       .io_requests_0_3_releaseLock( T2727 ),
       .io_requests_0_3_grant( swAllocator_io_requests_0_3_grant ),
       .io_requests_0_3_request( T2721 ),
       .io_requests_0_3_priorityLevel( R2717 ),
       .io_requests_0_2_releaseLock( T2713 ),
       .io_requests_0_2_grant( swAllocator_io_requests_0_2_grant ),
       .io_requests_0_2_request( T2707 ),
       .io_requests_0_2_priorityLevel( R2703 ),
       .io_requests_0_1_releaseLock( T2699 ),
       .io_requests_0_1_grant( swAllocator_io_requests_0_1_grant ),
       .io_requests_0_1_request( T2693 ),
       .io_requests_0_1_priorityLevel( R2689 ),
       .io_requests_0_0_releaseLock( T2685 ),
       .io_requests_0_0_grant( swAllocator_io_requests_0_0_grant ),
       .io_requests_0_0_request( T2679 ),
       .io_requests_0_0_priorityLevel( R2675 ),
       .io_resources_4_ready( 1'h1 ),
       //.io_resources_4_valid(  )
       .io_resources_3_ready( 1'h1 ),
       //.io_resources_3_valid(  )
       .io_resources_2_ready( 1'h1 ),
       //.io_resources_2_valid(  )
       .io_resources_1_ready( 1'h1 ),
       //.io_resources_1_valid(  )
       .io_resources_0_ready( 1'h1 ),
       //.io_resources_0_valid(  )
       .io_chosens_4( swAllocator_io_chosens_4 ),
       .io_chosens_3( swAllocator_io_chosens_3 ),
       .io_chosens_2( swAllocator_io_chosens_2 ),
       .io_chosens_1( swAllocator_io_chosens_1 ),
       .io_chosens_0( swAllocator_io_chosens_0 )
  );
  SwitchAllocator_1 vcAllocator(.clk(clk), .reset(reset),
       .io_requests_9_9_releaseLock( R2671 ),
       //.io_requests_9_9_grant(  )
       .io_requests_9_9_request( T2670 ),
       //.io_requests_9_9_priorityLevel(  )
       .io_requests_9_8_releaseLock( R2666 ),
       //.io_requests_9_8_grant(  )
       .io_requests_9_8_request( T2665 ),
       //.io_requests_9_8_priorityLevel(  )
       .io_requests_9_7_releaseLock( R2661 ),
       //.io_requests_9_7_grant(  )
       .io_requests_9_7_request( T2660 ),
       //.io_requests_9_7_priorityLevel(  )
       .io_requests_9_6_releaseLock( R2656 ),
       //.io_requests_9_6_grant(  )
       .io_requests_9_6_request( T2655 ),
       //.io_requests_9_6_priorityLevel(  )
       .io_requests_9_5_releaseLock( R2651 ),
       //.io_requests_9_5_grant(  )
       .io_requests_9_5_request( T2650 ),
       //.io_requests_9_5_priorityLevel(  )
       .io_requests_9_4_releaseLock( R2646 ),
       //.io_requests_9_4_grant(  )
       .io_requests_9_4_request( T2645 ),
       //.io_requests_9_4_priorityLevel(  )
       .io_requests_9_3_releaseLock( R2641 ),
       //.io_requests_9_3_grant(  )
       .io_requests_9_3_request( T2640 ),
       //.io_requests_9_3_priorityLevel(  )
       .io_requests_9_2_releaseLock( R2636 ),
       //.io_requests_9_2_grant(  )
       .io_requests_9_2_request( T2635 ),
       //.io_requests_9_2_priorityLevel(  )
       .io_requests_9_1_releaseLock( R2631 ),
       //.io_requests_9_1_grant(  )
       .io_requests_9_1_request( T2630 ),
       //.io_requests_9_1_priorityLevel(  )
       .io_requests_9_0_releaseLock( R2626 ),
       //.io_requests_9_0_grant(  )
       .io_requests_9_0_request( T2625 ),
       //.io_requests_9_0_priorityLevel(  )
       .io_requests_8_9_releaseLock( R2621 ),
       //.io_requests_8_9_grant(  )
       .io_requests_8_9_request( T2620 ),
       //.io_requests_8_9_priorityLevel(  )
       .io_requests_8_8_releaseLock( R2616 ),
       //.io_requests_8_8_grant(  )
       .io_requests_8_8_request( T2615 ),
       //.io_requests_8_8_priorityLevel(  )
       .io_requests_8_7_releaseLock( R2611 ),
       //.io_requests_8_7_grant(  )
       .io_requests_8_7_request( T2610 ),
       //.io_requests_8_7_priorityLevel(  )
       .io_requests_8_6_releaseLock( R2606 ),
       //.io_requests_8_6_grant(  )
       .io_requests_8_6_request( T2605 ),
       //.io_requests_8_6_priorityLevel(  )
       .io_requests_8_5_releaseLock( R2601 ),
       //.io_requests_8_5_grant(  )
       .io_requests_8_5_request( T2600 ),
       //.io_requests_8_5_priorityLevel(  )
       .io_requests_8_4_releaseLock( R2596 ),
       //.io_requests_8_4_grant(  )
       .io_requests_8_4_request( T2595 ),
       //.io_requests_8_4_priorityLevel(  )
       .io_requests_8_3_releaseLock( R2591 ),
       //.io_requests_8_3_grant(  )
       .io_requests_8_3_request( T2590 ),
       //.io_requests_8_3_priorityLevel(  )
       .io_requests_8_2_releaseLock( R2586 ),
       //.io_requests_8_2_grant(  )
       .io_requests_8_2_request( T2585 ),
       //.io_requests_8_2_priorityLevel(  )
       .io_requests_8_1_releaseLock( R2581 ),
       //.io_requests_8_1_grant(  )
       .io_requests_8_1_request( T2580 ),
       //.io_requests_8_1_priorityLevel(  )
       .io_requests_8_0_releaseLock( R2576 ),
       //.io_requests_8_0_grant(  )
       .io_requests_8_0_request( T2575 ),
       //.io_requests_8_0_priorityLevel(  )
       .io_requests_7_9_releaseLock( R2571 ),
       //.io_requests_7_9_grant(  )
       .io_requests_7_9_request( T2570 ),
       //.io_requests_7_9_priorityLevel(  )
       .io_requests_7_8_releaseLock( R2566 ),
       //.io_requests_7_8_grant(  )
       .io_requests_7_8_request( T2565 ),
       //.io_requests_7_8_priorityLevel(  )
       .io_requests_7_7_releaseLock( R2561 ),
       //.io_requests_7_7_grant(  )
       .io_requests_7_7_request( T2560 ),
       //.io_requests_7_7_priorityLevel(  )
       .io_requests_7_6_releaseLock( R2556 ),
       //.io_requests_7_6_grant(  )
       .io_requests_7_6_request( T2555 ),
       //.io_requests_7_6_priorityLevel(  )
       .io_requests_7_5_releaseLock( R2551 ),
       //.io_requests_7_5_grant(  )
       .io_requests_7_5_request( T2550 ),
       //.io_requests_7_5_priorityLevel(  )
       .io_requests_7_4_releaseLock( R2546 ),
       //.io_requests_7_4_grant(  )
       .io_requests_7_4_request( T2545 ),
       //.io_requests_7_4_priorityLevel(  )
       .io_requests_7_3_releaseLock( R2541 ),
       //.io_requests_7_3_grant(  )
       .io_requests_7_3_request( T2540 ),
       //.io_requests_7_3_priorityLevel(  )
       .io_requests_7_2_releaseLock( R2536 ),
       //.io_requests_7_2_grant(  )
       .io_requests_7_2_request( T2535 ),
       //.io_requests_7_2_priorityLevel(  )
       .io_requests_7_1_releaseLock( R2531 ),
       //.io_requests_7_1_grant(  )
       .io_requests_7_1_request( T2530 ),
       //.io_requests_7_1_priorityLevel(  )
       .io_requests_7_0_releaseLock( R2526 ),
       //.io_requests_7_0_grant(  )
       .io_requests_7_0_request( T2525 ),
       //.io_requests_7_0_priorityLevel(  )
       .io_requests_6_9_releaseLock( R2521 ),
       //.io_requests_6_9_grant(  )
       .io_requests_6_9_request( T2520 ),
       //.io_requests_6_9_priorityLevel(  )
       .io_requests_6_8_releaseLock( R2516 ),
       //.io_requests_6_8_grant(  )
       .io_requests_6_8_request( T2515 ),
       //.io_requests_6_8_priorityLevel(  )
       .io_requests_6_7_releaseLock( R2511 ),
       //.io_requests_6_7_grant(  )
       .io_requests_6_7_request( T2510 ),
       //.io_requests_6_7_priorityLevel(  )
       .io_requests_6_6_releaseLock( R2506 ),
       //.io_requests_6_6_grant(  )
       .io_requests_6_6_request( T2505 ),
       //.io_requests_6_6_priorityLevel(  )
       .io_requests_6_5_releaseLock( R2501 ),
       //.io_requests_6_5_grant(  )
       .io_requests_6_5_request( T2500 ),
       //.io_requests_6_5_priorityLevel(  )
       .io_requests_6_4_releaseLock( R2496 ),
       //.io_requests_6_4_grant(  )
       .io_requests_6_4_request( T2495 ),
       //.io_requests_6_4_priorityLevel(  )
       .io_requests_6_3_releaseLock( R2491 ),
       //.io_requests_6_3_grant(  )
       .io_requests_6_3_request( T2490 ),
       //.io_requests_6_3_priorityLevel(  )
       .io_requests_6_2_releaseLock( R2486 ),
       //.io_requests_6_2_grant(  )
       .io_requests_6_2_request( T2485 ),
       //.io_requests_6_2_priorityLevel(  )
       .io_requests_6_1_releaseLock( R2481 ),
       //.io_requests_6_1_grant(  )
       .io_requests_6_1_request( T2480 ),
       //.io_requests_6_1_priorityLevel(  )
       .io_requests_6_0_releaseLock( R2476 ),
       //.io_requests_6_0_grant(  )
       .io_requests_6_0_request( T2475 ),
       //.io_requests_6_0_priorityLevel(  )
       .io_requests_5_9_releaseLock( R2471 ),
       //.io_requests_5_9_grant(  )
       .io_requests_5_9_request( T2470 ),
       //.io_requests_5_9_priorityLevel(  )
       .io_requests_5_8_releaseLock( R2466 ),
       //.io_requests_5_8_grant(  )
       .io_requests_5_8_request( T2465 ),
       //.io_requests_5_8_priorityLevel(  )
       .io_requests_5_7_releaseLock( R2461 ),
       //.io_requests_5_7_grant(  )
       .io_requests_5_7_request( T2460 ),
       //.io_requests_5_7_priorityLevel(  )
       .io_requests_5_6_releaseLock( R2456 ),
       //.io_requests_5_6_grant(  )
       .io_requests_5_6_request( T2455 ),
       //.io_requests_5_6_priorityLevel(  )
       .io_requests_5_5_releaseLock( R2451 ),
       //.io_requests_5_5_grant(  )
       .io_requests_5_5_request( T2450 ),
       //.io_requests_5_5_priorityLevel(  )
       .io_requests_5_4_releaseLock( R2446 ),
       //.io_requests_5_4_grant(  )
       .io_requests_5_4_request( T2445 ),
       //.io_requests_5_4_priorityLevel(  )
       .io_requests_5_3_releaseLock( R2441 ),
       //.io_requests_5_3_grant(  )
       .io_requests_5_3_request( T2440 ),
       //.io_requests_5_3_priorityLevel(  )
       .io_requests_5_2_releaseLock( R2436 ),
       //.io_requests_5_2_grant(  )
       .io_requests_5_2_request( T2435 ),
       //.io_requests_5_2_priorityLevel(  )
       .io_requests_5_1_releaseLock( R2431 ),
       //.io_requests_5_1_grant(  )
       .io_requests_5_1_request( T2430 ),
       //.io_requests_5_1_priorityLevel(  )
       .io_requests_5_0_releaseLock( R2426 ),
       //.io_requests_5_0_grant(  )
       .io_requests_5_0_request( T2425 ),
       //.io_requests_5_0_priorityLevel(  )
       .io_requests_4_9_releaseLock( R2421 ),
       //.io_requests_4_9_grant(  )
       .io_requests_4_9_request( T2420 ),
       //.io_requests_4_9_priorityLevel(  )
       .io_requests_4_8_releaseLock( R2416 ),
       //.io_requests_4_8_grant(  )
       .io_requests_4_8_request( T2415 ),
       //.io_requests_4_8_priorityLevel(  )
       .io_requests_4_7_releaseLock( R2411 ),
       //.io_requests_4_7_grant(  )
       .io_requests_4_7_request( T2410 ),
       //.io_requests_4_7_priorityLevel(  )
       .io_requests_4_6_releaseLock( R2406 ),
       //.io_requests_4_6_grant(  )
       .io_requests_4_6_request( T2405 ),
       //.io_requests_4_6_priorityLevel(  )
       .io_requests_4_5_releaseLock( R2401 ),
       //.io_requests_4_5_grant(  )
       .io_requests_4_5_request( T2400 ),
       //.io_requests_4_5_priorityLevel(  )
       .io_requests_4_4_releaseLock( R2396 ),
       //.io_requests_4_4_grant(  )
       .io_requests_4_4_request( T2395 ),
       //.io_requests_4_4_priorityLevel(  )
       .io_requests_4_3_releaseLock( R2391 ),
       //.io_requests_4_3_grant(  )
       .io_requests_4_3_request( T2390 ),
       //.io_requests_4_3_priorityLevel(  )
       .io_requests_4_2_releaseLock( R2386 ),
       //.io_requests_4_2_grant(  )
       .io_requests_4_2_request( T2385 ),
       //.io_requests_4_2_priorityLevel(  )
       .io_requests_4_1_releaseLock( R2381 ),
       //.io_requests_4_1_grant(  )
       .io_requests_4_1_request( T2380 ),
       //.io_requests_4_1_priorityLevel(  )
       .io_requests_4_0_releaseLock( R2376 ),
       //.io_requests_4_0_grant(  )
       .io_requests_4_0_request( T2375 ),
       //.io_requests_4_0_priorityLevel(  )
       .io_requests_3_9_releaseLock( R2371 ),
       //.io_requests_3_9_grant(  )
       .io_requests_3_9_request( T2370 ),
       //.io_requests_3_9_priorityLevel(  )
       .io_requests_3_8_releaseLock( R2366 ),
       //.io_requests_3_8_grant(  )
       .io_requests_3_8_request( T2365 ),
       //.io_requests_3_8_priorityLevel(  )
       .io_requests_3_7_releaseLock( R2361 ),
       //.io_requests_3_7_grant(  )
       .io_requests_3_7_request( T2360 ),
       //.io_requests_3_7_priorityLevel(  )
       .io_requests_3_6_releaseLock( R2356 ),
       //.io_requests_3_6_grant(  )
       .io_requests_3_6_request( T2355 ),
       //.io_requests_3_6_priorityLevel(  )
       .io_requests_3_5_releaseLock( R2351 ),
       //.io_requests_3_5_grant(  )
       .io_requests_3_5_request( T2350 ),
       //.io_requests_3_5_priorityLevel(  )
       .io_requests_3_4_releaseLock( R2346 ),
       //.io_requests_3_4_grant(  )
       .io_requests_3_4_request( T2345 ),
       //.io_requests_3_4_priorityLevel(  )
       .io_requests_3_3_releaseLock( R2341 ),
       //.io_requests_3_3_grant(  )
       .io_requests_3_3_request( T2340 ),
       //.io_requests_3_3_priorityLevel(  )
       .io_requests_3_2_releaseLock( R2336 ),
       //.io_requests_3_2_grant(  )
       .io_requests_3_2_request( T2335 ),
       //.io_requests_3_2_priorityLevel(  )
       .io_requests_3_1_releaseLock( R2331 ),
       //.io_requests_3_1_grant(  )
       .io_requests_3_1_request( T2330 ),
       //.io_requests_3_1_priorityLevel(  )
       .io_requests_3_0_releaseLock( R2326 ),
       //.io_requests_3_0_grant(  )
       .io_requests_3_0_request( T2325 ),
       //.io_requests_3_0_priorityLevel(  )
       .io_requests_2_9_releaseLock( R2321 ),
       //.io_requests_2_9_grant(  )
       .io_requests_2_9_request( T2320 ),
       //.io_requests_2_9_priorityLevel(  )
       .io_requests_2_8_releaseLock( R2316 ),
       //.io_requests_2_8_grant(  )
       .io_requests_2_8_request( T2315 ),
       //.io_requests_2_8_priorityLevel(  )
       .io_requests_2_7_releaseLock( R2311 ),
       //.io_requests_2_7_grant(  )
       .io_requests_2_7_request( T2310 ),
       //.io_requests_2_7_priorityLevel(  )
       .io_requests_2_6_releaseLock( R2306 ),
       //.io_requests_2_6_grant(  )
       .io_requests_2_6_request( T2305 ),
       //.io_requests_2_6_priorityLevel(  )
       .io_requests_2_5_releaseLock( R2301 ),
       //.io_requests_2_5_grant(  )
       .io_requests_2_5_request( T2300 ),
       //.io_requests_2_5_priorityLevel(  )
       .io_requests_2_4_releaseLock( R2296 ),
       //.io_requests_2_4_grant(  )
       .io_requests_2_4_request( T2295 ),
       //.io_requests_2_4_priorityLevel(  )
       .io_requests_2_3_releaseLock( R2291 ),
       //.io_requests_2_3_grant(  )
       .io_requests_2_3_request( T2290 ),
       //.io_requests_2_3_priorityLevel(  )
       .io_requests_2_2_releaseLock( R2286 ),
       //.io_requests_2_2_grant(  )
       .io_requests_2_2_request( T2285 ),
       //.io_requests_2_2_priorityLevel(  )
       .io_requests_2_1_releaseLock( R2281 ),
       //.io_requests_2_1_grant(  )
       .io_requests_2_1_request( T2280 ),
       //.io_requests_2_1_priorityLevel(  )
       .io_requests_2_0_releaseLock( R2276 ),
       //.io_requests_2_0_grant(  )
       .io_requests_2_0_request( T2275 ),
       //.io_requests_2_0_priorityLevel(  )
       .io_requests_1_9_releaseLock( R2271 ),
       //.io_requests_1_9_grant(  )
       .io_requests_1_9_request( T2270 ),
       //.io_requests_1_9_priorityLevel(  )
       .io_requests_1_8_releaseLock( R2266 ),
       //.io_requests_1_8_grant(  )
       .io_requests_1_8_request( T2265 ),
       //.io_requests_1_8_priorityLevel(  )
       .io_requests_1_7_releaseLock( R2261 ),
       //.io_requests_1_7_grant(  )
       .io_requests_1_7_request( T2260 ),
       //.io_requests_1_7_priorityLevel(  )
       .io_requests_1_6_releaseLock( R2256 ),
       //.io_requests_1_6_grant(  )
       .io_requests_1_6_request( T2255 ),
       //.io_requests_1_6_priorityLevel(  )
       .io_requests_1_5_releaseLock( R2251 ),
       //.io_requests_1_5_grant(  )
       .io_requests_1_5_request( T2250 ),
       //.io_requests_1_5_priorityLevel(  )
       .io_requests_1_4_releaseLock( R2246 ),
       //.io_requests_1_4_grant(  )
       .io_requests_1_4_request( T2245 ),
       //.io_requests_1_4_priorityLevel(  )
       .io_requests_1_3_releaseLock( R2241 ),
       //.io_requests_1_3_grant(  )
       .io_requests_1_3_request( T2240 ),
       //.io_requests_1_3_priorityLevel(  )
       .io_requests_1_2_releaseLock( R2236 ),
       //.io_requests_1_2_grant(  )
       .io_requests_1_2_request( T2235 ),
       //.io_requests_1_2_priorityLevel(  )
       .io_requests_1_1_releaseLock( R2231 ),
       //.io_requests_1_1_grant(  )
       .io_requests_1_1_request( T2230 ),
       //.io_requests_1_1_priorityLevel(  )
       .io_requests_1_0_releaseLock( R2226 ),
       //.io_requests_1_0_grant(  )
       .io_requests_1_0_request( T2225 ),
       //.io_requests_1_0_priorityLevel(  )
       .io_requests_0_9_releaseLock( R2221 ),
       //.io_requests_0_9_grant(  )
       .io_requests_0_9_request( T2220 ),
       //.io_requests_0_9_priorityLevel(  )
       .io_requests_0_8_releaseLock( R2216 ),
       //.io_requests_0_8_grant(  )
       .io_requests_0_8_request( T2215 ),
       //.io_requests_0_8_priorityLevel(  )
       .io_requests_0_7_releaseLock( R2211 ),
       //.io_requests_0_7_grant(  )
       .io_requests_0_7_request( T2210 ),
       //.io_requests_0_7_priorityLevel(  )
       .io_requests_0_6_releaseLock( R2206 ),
       //.io_requests_0_6_grant(  )
       .io_requests_0_6_request( T2205 ),
       //.io_requests_0_6_priorityLevel(  )
       .io_requests_0_5_releaseLock( R2201 ),
       //.io_requests_0_5_grant(  )
       .io_requests_0_5_request( T2200 ),
       //.io_requests_0_5_priorityLevel(  )
       .io_requests_0_4_releaseLock( R2196 ),
       //.io_requests_0_4_grant(  )
       .io_requests_0_4_request( T2195 ),
       //.io_requests_0_4_priorityLevel(  )
       .io_requests_0_3_releaseLock( R2191 ),
       //.io_requests_0_3_grant(  )
       .io_requests_0_3_request( T2190 ),
       //.io_requests_0_3_priorityLevel(  )
       .io_requests_0_2_releaseLock( R2186 ),
       //.io_requests_0_2_grant(  )
       .io_requests_0_2_request( T2185 ),
       //.io_requests_0_2_priorityLevel(  )
       .io_requests_0_1_releaseLock( R2181 ),
       //.io_requests_0_1_grant(  )
       .io_requests_0_1_request( T2180 ),
       //.io_requests_0_1_priorityLevel(  )
       .io_requests_0_0_releaseLock( R2176 ),
       //.io_requests_0_0_grant(  )
       .io_requests_0_0_request( T2175 ),
       //.io_requests_0_0_priorityLevel(  )
       .io_resources_9_ready( T2173 ),
       .io_resources_9_valid( vcAllocator_io_resources_9_valid ),
       .io_resources_8_ready( T2171 ),
       .io_resources_8_valid( vcAllocator_io_resources_8_valid ),
       .io_resources_7_ready( T2169 ),
       .io_resources_7_valid( vcAllocator_io_resources_7_valid ),
       .io_resources_6_ready( T2167 ),
       .io_resources_6_valid( vcAllocator_io_resources_6_valid ),
       .io_resources_5_ready( T2165 ),
       .io_resources_5_valid( vcAllocator_io_resources_5_valid ),
       .io_resources_4_ready( T2163 ),
       .io_resources_4_valid( vcAllocator_io_resources_4_valid ),
       .io_resources_3_ready( T2161 ),
       .io_resources_3_valid( vcAllocator_io_resources_3_valid ),
       .io_resources_2_ready( T2159 ),
       .io_resources_2_valid( vcAllocator_io_resources_2_valid ),
       .io_resources_1_ready( T2157 ),
       .io_resources_1_valid( vcAllocator_io_resources_1_valid ),
       .io_resources_0_ready( T2155 ),
       .io_resources_0_valid( vcAllocator_io_resources_0_valid ),
       .io_chosens_9( vcAllocator_io_chosens_9 ),
       .io_chosens_8( vcAllocator_io_chosens_8 ),
       .io_chosens_7( vcAllocator_io_chosens_7 ),
       .io_chosens_6( vcAllocator_io_chosens_6 ),
       .io_chosens_5( vcAllocator_io_chosens_5 ),
       .io_chosens_4( vcAllocator_io_chosens_4 ),
       .io_chosens_3( vcAllocator_io_chosens_3 ),
       .io_chosens_2( vcAllocator_io_chosens_2 ),
       .io_chosens_1( vcAllocator_io_chosens_1 ),
       .io_chosens_0( vcAllocator_io_chosens_0 )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign vcAllocator.io_requests_9_9_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_9_8_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_9_7_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_9_6_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_9_5_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_9_4_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_9_3_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_9_2_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_9_1_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_9_0_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_8_9_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_8_8_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_8_7_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_8_6_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_8_5_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_8_4_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_8_3_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_8_2_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_8_1_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_8_0_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_7_9_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_7_8_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_7_7_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_7_6_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_7_5_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_7_4_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_7_3_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_7_2_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_7_1_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_7_0_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_6_9_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_6_8_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_6_7_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_6_6_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_6_5_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_6_4_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_6_3_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_6_2_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_6_1_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_6_0_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_5_9_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_5_8_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_5_7_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_5_6_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_5_5_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_5_4_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_5_3_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_5_2_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_5_1_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_5_0_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_4_9_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_4_8_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_4_7_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_4_6_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_4_5_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_4_4_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_4_3_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_4_2_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_4_1_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_4_0_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_3_9_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_3_8_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_3_7_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_3_6_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_3_5_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_3_4_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_3_3_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_3_2_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_3_1_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_3_0_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_2_9_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_2_8_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_2_7_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_2_6_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_2_5_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_2_4_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_2_3_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_2_2_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_2_1_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_2_0_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_1_9_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_1_8_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_1_7_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_1_6_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_1_5_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_1_4_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_1_3_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_1_2_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_1_1_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_1_0_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_0_9_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_0_8_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_0_7_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_0_6_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_0_5_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_0_4_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_0_3_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_0_2_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_0_1_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_0_0_priorityLevel = {1{1'b0}};
// synthesis translate_on
`endif
  VCRouterOutputStateManagement VCRouterOutputStateManagement(.clk(clk), .reset(reset),
       .io_swAllocGranted( T2094 ),
       .io_creditsAvail( T2092 ),
       .io_currentState( VCRouterOutputStateManagement_io_currentState )
  );
  VCRouterOutputStateManagement VCRouterOutputStateManagement_1(.clk(clk), .reset(reset),
       .io_swAllocGranted( T2031 ),
       .io_creditsAvail( T2029 ),
       .io_currentState( VCRouterOutputStateManagement_1_io_currentState )
  );
  VCRouterOutputStateManagement VCRouterOutputStateManagement_2(.clk(clk), .reset(reset),
       .io_swAllocGranted( T1968 ),
       .io_creditsAvail( T1966 ),
       .io_currentState( VCRouterOutputStateManagement_2_io_currentState )
  );
  VCRouterOutputStateManagement VCRouterOutputStateManagement_3(.clk(clk), .reset(reset),
       .io_swAllocGranted( T1905 ),
       .io_creditsAvail( T1903 ),
       .io_currentState( VCRouterOutputStateManagement_3_io_currentState )
  );
  VCRouterOutputStateManagement VCRouterOutputStateManagement_4(.clk(clk), .reset(reset),
       .io_swAllocGranted( T1722 ),
       .io_creditsAvail( T1720 ),
       .io_currentState( VCRouterOutputStateManagement_4_io_currentState )
  );
  CreditGen CreditGen(
       .io_outCredit_grant( CreditGen_io_outCredit_grant ),
       .io_inGrant( T1710 )
  );
  RouterRegFile RouterRegFile(.clk(clk), .reset(reset),
       .io_writeData( T1708 ),
       .io_writeEnable( T1705 ),
       //.io_full(  )
       .io_readData( RouterRegFile_io_readData ),
       .io_readValid( RouterRegFile_io_readValid ),
       .io_readIncrement( T1692 ),
       .io_writePipelineReg_2( RouterRegFile_io_readPipelineReg_1 ),
       .io_writePipelineReg_1( RouterRegFile_io_readPipelineReg_0 ),
       .io_writePipelineReg_0( T3181 ),
       .io_wePipelineReg_2( T1681 ),
       .io_wePipelineReg_1( T1678 ),
       .io_wePipelineReg_0( T1676 ),
       //.io_readPipelineReg_2(  )
       .io_readPipelineReg_1( RouterRegFile_io_readPipelineReg_1 ),
       .io_readPipelineReg_0( RouterRegFile_io_readPipelineReg_0 ),
       //.io_rvPipelineReg_2(  )
       .io_rvPipelineReg_1( RouterRegFile_io_rvPipelineReg_1 ),
       .io_rvPipelineReg_0( RouterRegFile_io_rvPipelineReg_0 )
  );
  RouterBuffer RouterBuffer(.clk(clk), .reset(reset),
       .io_enq_ready( RouterBuffer_io_enq_ready ),
       .io_enq_valid( T1675 ),
       .io_enq_bits_x( io_inChannels_0_flit_x ),
       .io_deq_ready( T1656 ),
       .io_deq_valid( RouterBuffer_io_deq_valid ),
       .io_deq_bits_x( RouterBuffer_io_deq_bits_x )
  );
  CMeshDOR_1 CMeshDOR(
       .io_inHeadFlit_packetID( T1655 ),
       .io_inHeadFlit_isTail( T1654 ),
       .io_inHeadFlit_vcPort( T1653 ),
       .io_inHeadFlit_packetType( T1652 ),
       .io_inHeadFlit_destination_2( T1651 ),
       .io_inHeadFlit_destination_1( T1650 ),
       .io_inHeadFlit_destination_0( T1649 ),
       .io_inHeadFlit_priorityLevel( T1646 ),
       .io_outHeadFlit_packetID( CMeshDOR_io_outHeadFlit_packetID ),
       .io_outHeadFlit_isTail( CMeshDOR_io_outHeadFlit_isTail ),
       .io_outHeadFlit_vcPort( CMeshDOR_io_outHeadFlit_vcPort ),
       .io_outHeadFlit_packetType( CMeshDOR_io_outHeadFlit_packetType ),
       .io_outHeadFlit_destination_2( CMeshDOR_io_outHeadFlit_destination_2 ),
       .io_outHeadFlit_destination_1( CMeshDOR_io_outHeadFlit_destination_1 ),
       .io_outHeadFlit_destination_0( CMeshDOR_io_outHeadFlit_destination_0 ),
       .io_outHeadFlit_priorityLevel( CMeshDOR_io_outHeadFlit_priorityLevel ),
       .io_result( CMeshDOR_io_result ),
       .io_vcsAvailable_4( CMeshDOR_io_vcsAvailable_4 ),
       .io_vcsAvailable_3( CMeshDOR_io_vcsAvailable_3 ),
       .io_vcsAvailable_2( CMeshDOR_io_vcsAvailable_2 ),
       .io_vcsAvailable_1( CMeshDOR_io_vcsAvailable_1 ),
       .io_vcsAvailable_0( CMeshDOR_io_vcsAvailable_0 )
  );
  VCRouterStateManagement VCRouterStateManagement(.clk(clk), .reset(reset),
       .io_inputBufferValid( RouterBuffer_io_deq_valid ),
       .io_routingComplete( R1645 ),
       .io_inputBufferIsTail( T1636 ),
       .io_vcAllocGranted( vcAllocator_io_resources_0_valid ),
       .io_swAllocGranted( T1616 ),
       .io_creditsAvail( T1597 ),
       .io_outputReady( T1584 ),
       .io_currentState( VCRouterStateManagement_io_currentState )
  );
  ReplaceVCPort ReplaceVCPort(
       .io_oldFlit_x( T1582 ),
       .io_newVCPort( T3175 ),
       .io_newFlit_x( ReplaceVCPort_io_newFlit_x )
  );
  Flit2FlitBundle Flit2FlitBundle(
       .io_inFlit_x( T1576 )
       //.io_outHead_packetID(  )
       //.io_outHead_isTail(  )
       //.io_outHead_vcPort(  )
       //.io_outHead_packetType(  )
       //.io_outHead_destination_2(  )
       //.io_outHead_destination_1(  )
       //.io_outHead_destination_0(  )
       //.io_outHead_priorityLevel(  )
       //.io_outBody_packetID(  )
       //.io_outBody_isTail(  )
       //.io_outBody_vcPort(  )
       //.io_outBody_flitID(  )
       //.io_outBody_payload(  )
  );
  CreditGen CreditGen_1(
       .io_outCredit_grant( CreditGen_1_io_outCredit_grant ),
       .io_inGrant( T1566 )
  );
  RouterRegFile RouterRegFile_1(.clk(clk), .reset(reset),
       .io_writeData( T1564 ),
       .io_writeEnable( T1561 ),
       //.io_full(  )
       .io_readData( RouterRegFile_1_io_readData ),
       .io_readValid( RouterRegFile_1_io_readValid ),
       .io_readIncrement( T1548 ),
       .io_writePipelineReg_2( RouterRegFile_1_io_readPipelineReg_1 ),
       .io_writePipelineReg_1( RouterRegFile_1_io_readPipelineReg_0 ),
       .io_writePipelineReg_0( T3174 ),
       .io_wePipelineReg_2( T1537 ),
       .io_wePipelineReg_1( T1534 ),
       .io_wePipelineReg_0( T1532 ),
       //.io_readPipelineReg_2(  )
       .io_readPipelineReg_1( RouterRegFile_1_io_readPipelineReg_1 ),
       .io_readPipelineReg_0( RouterRegFile_1_io_readPipelineReg_0 ),
       //.io_rvPipelineReg_2(  )
       .io_rvPipelineReg_1( RouterRegFile_1_io_rvPipelineReg_1 ),
       .io_rvPipelineReg_0( RouterRegFile_1_io_rvPipelineReg_0 )
  );
  RouterBuffer RouterBuffer_1(.clk(clk), .reset(reset),
       .io_enq_ready( RouterBuffer_1_io_enq_ready ),
       .io_enq_valid( T1531 ),
       .io_enq_bits_x( io_inChannels_0_flit_x ),
       .io_deq_ready( T1512 ),
       .io_deq_valid( RouterBuffer_1_io_deq_valid ),
       .io_deq_bits_x( RouterBuffer_1_io_deq_bits_x )
  );
  CMeshDOR_1 CMeshDOR_1(
       .io_inHeadFlit_packetID( T1511 ),
       .io_inHeadFlit_isTail( T1510 ),
       .io_inHeadFlit_vcPort( T1509 ),
       .io_inHeadFlit_packetType( T1508 ),
       .io_inHeadFlit_destination_2( T1507 ),
       .io_inHeadFlit_destination_1( T1506 ),
       .io_inHeadFlit_destination_0( T1505 ),
       .io_inHeadFlit_priorityLevel( T1502 ),
       .io_outHeadFlit_packetID( CMeshDOR_1_io_outHeadFlit_packetID ),
       .io_outHeadFlit_isTail( CMeshDOR_1_io_outHeadFlit_isTail ),
       .io_outHeadFlit_vcPort( CMeshDOR_1_io_outHeadFlit_vcPort ),
       .io_outHeadFlit_packetType( CMeshDOR_1_io_outHeadFlit_packetType ),
       .io_outHeadFlit_destination_2( CMeshDOR_1_io_outHeadFlit_destination_2 ),
       .io_outHeadFlit_destination_1( CMeshDOR_1_io_outHeadFlit_destination_1 ),
       .io_outHeadFlit_destination_0( CMeshDOR_1_io_outHeadFlit_destination_0 ),
       .io_outHeadFlit_priorityLevel( CMeshDOR_1_io_outHeadFlit_priorityLevel ),
       .io_result( CMeshDOR_1_io_result ),
       .io_vcsAvailable_4( CMeshDOR_1_io_vcsAvailable_4 ),
       .io_vcsAvailable_3( CMeshDOR_1_io_vcsAvailable_3 ),
       .io_vcsAvailable_2( CMeshDOR_1_io_vcsAvailable_2 ),
       .io_vcsAvailable_1( CMeshDOR_1_io_vcsAvailable_1 ),
       .io_vcsAvailable_0( CMeshDOR_1_io_vcsAvailable_0 )
  );
  VCRouterStateManagement VCRouterStateManagement_1(.clk(clk), .reset(reset),
       .io_inputBufferValid( RouterBuffer_1_io_deq_valid ),
       .io_routingComplete( R1501 ),
       .io_inputBufferIsTail( T1492 ),
       .io_vcAllocGranted( vcAllocator_io_resources_1_valid ),
       .io_swAllocGranted( T1472 ),
       .io_creditsAvail( T1453 ),
       .io_outputReady( T1440 ),
       .io_currentState( VCRouterStateManagement_1_io_currentState )
  );
  ReplaceVCPort ReplaceVCPort_1(
       .io_oldFlit_x( T1438 ),
       .io_newVCPort( T3168 ),
       .io_newFlit_x( ReplaceVCPort_1_io_newFlit_x )
  );
  Flit2FlitBundle Flit2FlitBundle_1(
       .io_inFlit_x( T1432 )
       //.io_outHead_packetID(  )
       //.io_outHead_isTail(  )
       //.io_outHead_vcPort(  )
       //.io_outHead_packetType(  )
       //.io_outHead_destination_2(  )
       //.io_outHead_destination_1(  )
       //.io_outHead_destination_0(  )
       //.io_outHead_priorityLevel(  )
       //.io_outBody_packetID(  )
       //.io_outBody_isTail(  )
       //.io_outBody_vcPort(  )
       //.io_outBody_flitID(  )
       //.io_outBody_payload(  )
  );
  CreditGen CreditGen_2(
       .io_outCredit_grant( CreditGen_2_io_outCredit_grant ),
       .io_inGrant( T1422 )
  );
  RouterRegFile RouterRegFile_2(.clk(clk), .reset(reset),
       .io_writeData( T1420 ),
       .io_writeEnable( T1417 ),
       //.io_full(  )
       .io_readData( RouterRegFile_2_io_readData ),
       .io_readValid( RouterRegFile_2_io_readValid ),
       .io_readIncrement( T1404 ),
       .io_writePipelineReg_2( RouterRegFile_2_io_readPipelineReg_1 ),
       .io_writePipelineReg_1( RouterRegFile_2_io_readPipelineReg_0 ),
       .io_writePipelineReg_0( T3167 ),
       .io_wePipelineReg_2( T1393 ),
       .io_wePipelineReg_1( T1390 ),
       .io_wePipelineReg_0( T1388 ),
       //.io_readPipelineReg_2(  )
       .io_readPipelineReg_1( RouterRegFile_2_io_readPipelineReg_1 ),
       .io_readPipelineReg_0( RouterRegFile_2_io_readPipelineReg_0 ),
       //.io_rvPipelineReg_2(  )
       .io_rvPipelineReg_1( RouterRegFile_2_io_rvPipelineReg_1 ),
       .io_rvPipelineReg_0( RouterRegFile_2_io_rvPipelineReg_0 )
  );
  RouterBuffer RouterBuffer_2(.clk(clk), .reset(reset),
       .io_enq_ready( RouterBuffer_2_io_enq_ready ),
       .io_enq_valid( T1387 ),
       .io_enq_bits_x( io_inChannels_1_flit_x ),
       .io_deq_ready( T1368 ),
       .io_deq_valid( RouterBuffer_2_io_deq_valid ),
       .io_deq_bits_x( RouterBuffer_2_io_deq_bits_x )
  );
  CMeshDOR_1 CMeshDOR_2(
       .io_inHeadFlit_packetID( T1367 ),
       .io_inHeadFlit_isTail( T1366 ),
       .io_inHeadFlit_vcPort( T1365 ),
       .io_inHeadFlit_packetType( T1364 ),
       .io_inHeadFlit_destination_2( T1363 ),
       .io_inHeadFlit_destination_1( T1362 ),
       .io_inHeadFlit_destination_0( T1361 ),
       .io_inHeadFlit_priorityLevel( T1358 ),
       .io_outHeadFlit_packetID( CMeshDOR_2_io_outHeadFlit_packetID ),
       .io_outHeadFlit_isTail( CMeshDOR_2_io_outHeadFlit_isTail ),
       .io_outHeadFlit_vcPort( CMeshDOR_2_io_outHeadFlit_vcPort ),
       .io_outHeadFlit_packetType( CMeshDOR_2_io_outHeadFlit_packetType ),
       .io_outHeadFlit_destination_2( CMeshDOR_2_io_outHeadFlit_destination_2 ),
       .io_outHeadFlit_destination_1( CMeshDOR_2_io_outHeadFlit_destination_1 ),
       .io_outHeadFlit_destination_0( CMeshDOR_2_io_outHeadFlit_destination_0 ),
       .io_outHeadFlit_priorityLevel( CMeshDOR_2_io_outHeadFlit_priorityLevel ),
       .io_result( CMeshDOR_2_io_result ),
       .io_vcsAvailable_4( CMeshDOR_2_io_vcsAvailable_4 ),
       .io_vcsAvailable_3( CMeshDOR_2_io_vcsAvailable_3 ),
       .io_vcsAvailable_2( CMeshDOR_2_io_vcsAvailable_2 ),
       .io_vcsAvailable_1( CMeshDOR_2_io_vcsAvailable_1 ),
       .io_vcsAvailable_0( CMeshDOR_2_io_vcsAvailable_0 )
  );
  VCRouterStateManagement VCRouterStateManagement_2(.clk(clk), .reset(reset),
       .io_inputBufferValid( RouterBuffer_2_io_deq_valid ),
       .io_routingComplete( R1357 ),
       .io_inputBufferIsTail( T1348 ),
       .io_vcAllocGranted( vcAllocator_io_resources_2_valid ),
       .io_swAllocGranted( T1328 ),
       .io_creditsAvail( T1309 ),
       .io_outputReady( T1296 ),
       .io_currentState( VCRouterStateManagement_2_io_currentState )
  );
  ReplaceVCPort ReplaceVCPort_2(
       .io_oldFlit_x( T1294 ),
       .io_newVCPort( T3161 ),
       .io_newFlit_x( ReplaceVCPort_2_io_newFlit_x )
  );
  Flit2FlitBundle Flit2FlitBundle_2(
       .io_inFlit_x( T1288 )
       //.io_outHead_packetID(  )
       //.io_outHead_isTail(  )
       //.io_outHead_vcPort(  )
       //.io_outHead_packetType(  )
       //.io_outHead_destination_2(  )
       //.io_outHead_destination_1(  )
       //.io_outHead_destination_0(  )
       //.io_outHead_priorityLevel(  )
       //.io_outBody_packetID(  )
       //.io_outBody_isTail(  )
       //.io_outBody_vcPort(  )
       //.io_outBody_flitID(  )
       //.io_outBody_payload(  )
  );
  CreditGen CreditGen_3(
       .io_outCredit_grant( CreditGen_3_io_outCredit_grant ),
       .io_inGrant( T1278 )
  );
  RouterRegFile RouterRegFile_3(.clk(clk), .reset(reset),
       .io_writeData( T1276 ),
       .io_writeEnable( T1273 ),
       //.io_full(  )
       .io_readData( RouterRegFile_3_io_readData ),
       .io_readValid( RouterRegFile_3_io_readValid ),
       .io_readIncrement( T1260 ),
       .io_writePipelineReg_2( RouterRegFile_3_io_readPipelineReg_1 ),
       .io_writePipelineReg_1( RouterRegFile_3_io_readPipelineReg_0 ),
       .io_writePipelineReg_0( T3160 ),
       .io_wePipelineReg_2( T1249 ),
       .io_wePipelineReg_1( T1246 ),
       .io_wePipelineReg_0( T1244 ),
       //.io_readPipelineReg_2(  )
       .io_readPipelineReg_1( RouterRegFile_3_io_readPipelineReg_1 ),
       .io_readPipelineReg_0( RouterRegFile_3_io_readPipelineReg_0 ),
       //.io_rvPipelineReg_2(  )
       .io_rvPipelineReg_1( RouterRegFile_3_io_rvPipelineReg_1 ),
       .io_rvPipelineReg_0( RouterRegFile_3_io_rvPipelineReg_0 )
  );
  RouterBuffer RouterBuffer_3(.clk(clk), .reset(reset),
       .io_enq_ready( RouterBuffer_3_io_enq_ready ),
       .io_enq_valid( T1243 ),
       .io_enq_bits_x( io_inChannels_1_flit_x ),
       .io_deq_ready( T1224 ),
       .io_deq_valid( RouterBuffer_3_io_deq_valid ),
       .io_deq_bits_x( RouterBuffer_3_io_deq_bits_x )
  );
  CMeshDOR_1 CMeshDOR_3(
       .io_inHeadFlit_packetID( T1223 ),
       .io_inHeadFlit_isTail( T1222 ),
       .io_inHeadFlit_vcPort( T1221 ),
       .io_inHeadFlit_packetType( T1220 ),
       .io_inHeadFlit_destination_2( T1219 ),
       .io_inHeadFlit_destination_1( T1218 ),
       .io_inHeadFlit_destination_0( T1217 ),
       .io_inHeadFlit_priorityLevel( T1214 ),
       .io_outHeadFlit_packetID( CMeshDOR_3_io_outHeadFlit_packetID ),
       .io_outHeadFlit_isTail( CMeshDOR_3_io_outHeadFlit_isTail ),
       .io_outHeadFlit_vcPort( CMeshDOR_3_io_outHeadFlit_vcPort ),
       .io_outHeadFlit_packetType( CMeshDOR_3_io_outHeadFlit_packetType ),
       .io_outHeadFlit_destination_2( CMeshDOR_3_io_outHeadFlit_destination_2 ),
       .io_outHeadFlit_destination_1( CMeshDOR_3_io_outHeadFlit_destination_1 ),
       .io_outHeadFlit_destination_0( CMeshDOR_3_io_outHeadFlit_destination_0 ),
       .io_outHeadFlit_priorityLevel( CMeshDOR_3_io_outHeadFlit_priorityLevel ),
       .io_result( CMeshDOR_3_io_result ),
       .io_vcsAvailable_4( CMeshDOR_3_io_vcsAvailable_4 ),
       .io_vcsAvailable_3( CMeshDOR_3_io_vcsAvailable_3 ),
       .io_vcsAvailable_2( CMeshDOR_3_io_vcsAvailable_2 ),
       .io_vcsAvailable_1( CMeshDOR_3_io_vcsAvailable_1 ),
       .io_vcsAvailable_0( CMeshDOR_3_io_vcsAvailable_0 )
  );
  VCRouterStateManagement VCRouterStateManagement_3(.clk(clk), .reset(reset),
       .io_inputBufferValid( RouterBuffer_3_io_deq_valid ),
       .io_routingComplete( R1213 ),
       .io_inputBufferIsTail( T1204 ),
       .io_vcAllocGranted( vcAllocator_io_resources_3_valid ),
       .io_swAllocGranted( T1184 ),
       .io_creditsAvail( T1165 ),
       .io_outputReady( T1152 ),
       .io_currentState( VCRouterStateManagement_3_io_currentState )
  );
  ReplaceVCPort ReplaceVCPort_3(
       .io_oldFlit_x( T1150 ),
       .io_newVCPort( T3154 ),
       .io_newFlit_x( ReplaceVCPort_3_io_newFlit_x )
  );
  Flit2FlitBundle Flit2FlitBundle_3(
       .io_inFlit_x( T1144 )
       //.io_outHead_packetID(  )
       //.io_outHead_isTail(  )
       //.io_outHead_vcPort(  )
       //.io_outHead_packetType(  )
       //.io_outHead_destination_2(  )
       //.io_outHead_destination_1(  )
       //.io_outHead_destination_0(  )
       //.io_outHead_priorityLevel(  )
       //.io_outBody_packetID(  )
       //.io_outBody_isTail(  )
       //.io_outBody_vcPort(  )
       //.io_outBody_flitID(  )
       //.io_outBody_payload(  )
  );
  CreditGen CreditGen_4(
       .io_outCredit_grant( CreditGen_4_io_outCredit_grant ),
       .io_inGrant( T1134 )
  );
  RouterRegFile RouterRegFile_4(.clk(clk), .reset(reset),
       .io_writeData( T1132 ),
       .io_writeEnable( T1129 ),
       //.io_full(  )
       .io_readData( RouterRegFile_4_io_readData ),
       .io_readValid( RouterRegFile_4_io_readValid ),
       .io_readIncrement( T1116 ),
       .io_writePipelineReg_2( RouterRegFile_4_io_readPipelineReg_1 ),
       .io_writePipelineReg_1( RouterRegFile_4_io_readPipelineReg_0 ),
       .io_writePipelineReg_0( T3153 ),
       .io_wePipelineReg_2( T1105 ),
       .io_wePipelineReg_1( T1102 ),
       .io_wePipelineReg_0( T1100 ),
       //.io_readPipelineReg_2(  )
       .io_readPipelineReg_1( RouterRegFile_4_io_readPipelineReg_1 ),
       .io_readPipelineReg_0( RouterRegFile_4_io_readPipelineReg_0 ),
       //.io_rvPipelineReg_2(  )
       .io_rvPipelineReg_1( RouterRegFile_4_io_rvPipelineReg_1 ),
       .io_rvPipelineReg_0( RouterRegFile_4_io_rvPipelineReg_0 )
  );
  RouterBuffer RouterBuffer_4(.clk(clk), .reset(reset),
       .io_enq_ready( RouterBuffer_4_io_enq_ready ),
       .io_enq_valid( T1099 ),
       .io_enq_bits_x( io_inChannels_2_flit_x ),
       .io_deq_ready( T1080 ),
       .io_deq_valid( RouterBuffer_4_io_deq_valid ),
       .io_deq_bits_x( RouterBuffer_4_io_deq_bits_x )
  );
  CMeshDOR_1 CMeshDOR_4(
       .io_inHeadFlit_packetID( T1079 ),
       .io_inHeadFlit_isTail( T1078 ),
       .io_inHeadFlit_vcPort( T1077 ),
       .io_inHeadFlit_packetType( T1076 ),
       .io_inHeadFlit_destination_2( T1075 ),
       .io_inHeadFlit_destination_1( T1074 ),
       .io_inHeadFlit_destination_0( T1073 ),
       .io_inHeadFlit_priorityLevel( T1070 ),
       .io_outHeadFlit_packetID( CMeshDOR_4_io_outHeadFlit_packetID ),
       .io_outHeadFlit_isTail( CMeshDOR_4_io_outHeadFlit_isTail ),
       .io_outHeadFlit_vcPort( CMeshDOR_4_io_outHeadFlit_vcPort ),
       .io_outHeadFlit_packetType( CMeshDOR_4_io_outHeadFlit_packetType ),
       .io_outHeadFlit_destination_2( CMeshDOR_4_io_outHeadFlit_destination_2 ),
       .io_outHeadFlit_destination_1( CMeshDOR_4_io_outHeadFlit_destination_1 ),
       .io_outHeadFlit_destination_0( CMeshDOR_4_io_outHeadFlit_destination_0 ),
       .io_outHeadFlit_priorityLevel( CMeshDOR_4_io_outHeadFlit_priorityLevel ),
       .io_result( CMeshDOR_4_io_result ),
       .io_vcsAvailable_4( CMeshDOR_4_io_vcsAvailable_4 ),
       .io_vcsAvailable_3( CMeshDOR_4_io_vcsAvailable_3 ),
       .io_vcsAvailable_2( CMeshDOR_4_io_vcsAvailable_2 ),
       .io_vcsAvailable_1( CMeshDOR_4_io_vcsAvailable_1 ),
       .io_vcsAvailable_0( CMeshDOR_4_io_vcsAvailable_0 )
  );
  VCRouterStateManagement VCRouterStateManagement_4(.clk(clk), .reset(reset),
       .io_inputBufferValid( RouterBuffer_4_io_deq_valid ),
       .io_routingComplete( R1069 ),
       .io_inputBufferIsTail( T1060 ),
       .io_vcAllocGranted( vcAllocator_io_resources_4_valid ),
       .io_swAllocGranted( T1040 ),
       .io_creditsAvail( T1021 ),
       .io_outputReady( T1008 ),
       .io_currentState( VCRouterStateManagement_4_io_currentState )
  );
  ReplaceVCPort ReplaceVCPort_4(
       .io_oldFlit_x( T1006 ),
       .io_newVCPort( T3147 ),
       .io_newFlit_x( ReplaceVCPort_4_io_newFlit_x )
  );
  Flit2FlitBundle Flit2FlitBundle_4(
       .io_inFlit_x( T1000 )
       //.io_outHead_packetID(  )
       //.io_outHead_isTail(  )
       //.io_outHead_vcPort(  )
       //.io_outHead_packetType(  )
       //.io_outHead_destination_2(  )
       //.io_outHead_destination_1(  )
       //.io_outHead_destination_0(  )
       //.io_outHead_priorityLevel(  )
       //.io_outBody_packetID(  )
       //.io_outBody_isTail(  )
       //.io_outBody_vcPort(  )
       //.io_outBody_flitID(  )
       //.io_outBody_payload(  )
  );
  CreditGen CreditGen_5(
       .io_outCredit_grant( CreditGen_5_io_outCredit_grant ),
       .io_inGrant( T990 )
  );
  RouterRegFile RouterRegFile_5(.clk(clk), .reset(reset),
       .io_writeData( T988 ),
       .io_writeEnable( T985 ),
       //.io_full(  )
       .io_readData( RouterRegFile_5_io_readData ),
       .io_readValid( RouterRegFile_5_io_readValid ),
       .io_readIncrement( T972 ),
       .io_writePipelineReg_2( RouterRegFile_5_io_readPipelineReg_1 ),
       .io_writePipelineReg_1( RouterRegFile_5_io_readPipelineReg_0 ),
       .io_writePipelineReg_0( T3146 ),
       .io_wePipelineReg_2( T961 ),
       .io_wePipelineReg_1( T958 ),
       .io_wePipelineReg_0( T956 ),
       //.io_readPipelineReg_2(  )
       .io_readPipelineReg_1( RouterRegFile_5_io_readPipelineReg_1 ),
       .io_readPipelineReg_0( RouterRegFile_5_io_readPipelineReg_0 ),
       //.io_rvPipelineReg_2(  )
       .io_rvPipelineReg_1( RouterRegFile_5_io_rvPipelineReg_1 ),
       .io_rvPipelineReg_0( RouterRegFile_5_io_rvPipelineReg_0 )
  );
  RouterBuffer RouterBuffer_5(.clk(clk), .reset(reset),
       .io_enq_ready( RouterBuffer_5_io_enq_ready ),
       .io_enq_valid( T955 ),
       .io_enq_bits_x( io_inChannels_2_flit_x ),
       .io_deq_ready( T936 ),
       .io_deq_valid( RouterBuffer_5_io_deq_valid ),
       .io_deq_bits_x( RouterBuffer_5_io_deq_bits_x )
  );
  CMeshDOR_1 CMeshDOR_5(
       .io_inHeadFlit_packetID( T935 ),
       .io_inHeadFlit_isTail( T934 ),
       .io_inHeadFlit_vcPort( T933 ),
       .io_inHeadFlit_packetType( T932 ),
       .io_inHeadFlit_destination_2( T931 ),
       .io_inHeadFlit_destination_1( T930 ),
       .io_inHeadFlit_destination_0( T929 ),
       .io_inHeadFlit_priorityLevel( T926 ),
       .io_outHeadFlit_packetID( CMeshDOR_5_io_outHeadFlit_packetID ),
       .io_outHeadFlit_isTail( CMeshDOR_5_io_outHeadFlit_isTail ),
       .io_outHeadFlit_vcPort( CMeshDOR_5_io_outHeadFlit_vcPort ),
       .io_outHeadFlit_packetType( CMeshDOR_5_io_outHeadFlit_packetType ),
       .io_outHeadFlit_destination_2( CMeshDOR_5_io_outHeadFlit_destination_2 ),
       .io_outHeadFlit_destination_1( CMeshDOR_5_io_outHeadFlit_destination_1 ),
       .io_outHeadFlit_destination_0( CMeshDOR_5_io_outHeadFlit_destination_0 ),
       .io_outHeadFlit_priorityLevel( CMeshDOR_5_io_outHeadFlit_priorityLevel ),
       .io_result( CMeshDOR_5_io_result ),
       .io_vcsAvailable_4( CMeshDOR_5_io_vcsAvailable_4 ),
       .io_vcsAvailable_3( CMeshDOR_5_io_vcsAvailable_3 ),
       .io_vcsAvailable_2( CMeshDOR_5_io_vcsAvailable_2 ),
       .io_vcsAvailable_1( CMeshDOR_5_io_vcsAvailable_1 ),
       .io_vcsAvailable_0( CMeshDOR_5_io_vcsAvailable_0 )
  );
  VCRouterStateManagement VCRouterStateManagement_5(.clk(clk), .reset(reset),
       .io_inputBufferValid( RouterBuffer_5_io_deq_valid ),
       .io_routingComplete( R925 ),
       .io_inputBufferIsTail( T916 ),
       .io_vcAllocGranted( vcAllocator_io_resources_5_valid ),
       .io_swAllocGranted( T896 ),
       .io_creditsAvail( T877 ),
       .io_outputReady( T864 ),
       .io_currentState( VCRouterStateManagement_5_io_currentState )
  );
  ReplaceVCPort ReplaceVCPort_5(
       .io_oldFlit_x( T862 ),
       .io_newVCPort( T3140 ),
       .io_newFlit_x( ReplaceVCPort_5_io_newFlit_x )
  );
  Flit2FlitBundle Flit2FlitBundle_5(
       .io_inFlit_x( T856 )
       //.io_outHead_packetID(  )
       //.io_outHead_isTail(  )
       //.io_outHead_vcPort(  )
       //.io_outHead_packetType(  )
       //.io_outHead_destination_2(  )
       //.io_outHead_destination_1(  )
       //.io_outHead_destination_0(  )
       //.io_outHead_priorityLevel(  )
       //.io_outBody_packetID(  )
       //.io_outBody_isTail(  )
       //.io_outBody_vcPort(  )
       //.io_outBody_flitID(  )
       //.io_outBody_payload(  )
  );
  CreditGen CreditGen_6(
       .io_outCredit_grant( CreditGen_6_io_outCredit_grant ),
       .io_inGrant( T846 )
  );
  RouterRegFile RouterRegFile_6(.clk(clk), .reset(reset),
       .io_writeData( T844 ),
       .io_writeEnable( T841 ),
       //.io_full(  )
       .io_readData( RouterRegFile_6_io_readData ),
       .io_readValid( RouterRegFile_6_io_readValid ),
       .io_readIncrement( T828 ),
       .io_writePipelineReg_2( RouterRegFile_6_io_readPipelineReg_1 ),
       .io_writePipelineReg_1( RouterRegFile_6_io_readPipelineReg_0 ),
       .io_writePipelineReg_0( T3139 ),
       .io_wePipelineReg_2( T817 ),
       .io_wePipelineReg_1( T814 ),
       .io_wePipelineReg_0( T812 ),
       //.io_readPipelineReg_2(  )
       .io_readPipelineReg_1( RouterRegFile_6_io_readPipelineReg_1 ),
       .io_readPipelineReg_0( RouterRegFile_6_io_readPipelineReg_0 ),
       //.io_rvPipelineReg_2(  )
       .io_rvPipelineReg_1( RouterRegFile_6_io_rvPipelineReg_1 ),
       .io_rvPipelineReg_0( RouterRegFile_6_io_rvPipelineReg_0 )
  );
  RouterBuffer RouterBuffer_6(.clk(clk), .reset(reset),
       .io_enq_ready( RouterBuffer_6_io_enq_ready ),
       .io_enq_valid( T811 ),
       .io_enq_bits_x( io_inChannels_3_flit_x ),
       .io_deq_ready( T792 ),
       .io_deq_valid( RouterBuffer_6_io_deq_valid ),
       .io_deq_bits_x( RouterBuffer_6_io_deq_bits_x )
  );
  CMeshDOR_1 CMeshDOR_6(
       .io_inHeadFlit_packetID( T791 ),
       .io_inHeadFlit_isTail( T790 ),
       .io_inHeadFlit_vcPort( T789 ),
       .io_inHeadFlit_packetType( T788 ),
       .io_inHeadFlit_destination_2( T787 ),
       .io_inHeadFlit_destination_1( T786 ),
       .io_inHeadFlit_destination_0( T785 ),
       .io_inHeadFlit_priorityLevel( T782 ),
       .io_outHeadFlit_packetID( CMeshDOR_6_io_outHeadFlit_packetID ),
       .io_outHeadFlit_isTail( CMeshDOR_6_io_outHeadFlit_isTail ),
       .io_outHeadFlit_vcPort( CMeshDOR_6_io_outHeadFlit_vcPort ),
       .io_outHeadFlit_packetType( CMeshDOR_6_io_outHeadFlit_packetType ),
       .io_outHeadFlit_destination_2( CMeshDOR_6_io_outHeadFlit_destination_2 ),
       .io_outHeadFlit_destination_1( CMeshDOR_6_io_outHeadFlit_destination_1 ),
       .io_outHeadFlit_destination_0( CMeshDOR_6_io_outHeadFlit_destination_0 ),
       .io_outHeadFlit_priorityLevel( CMeshDOR_6_io_outHeadFlit_priorityLevel ),
       .io_result( CMeshDOR_6_io_result ),
       .io_vcsAvailable_4( CMeshDOR_6_io_vcsAvailable_4 ),
       .io_vcsAvailable_3( CMeshDOR_6_io_vcsAvailable_3 ),
       .io_vcsAvailable_2( CMeshDOR_6_io_vcsAvailable_2 ),
       .io_vcsAvailable_1( CMeshDOR_6_io_vcsAvailable_1 ),
       .io_vcsAvailable_0( CMeshDOR_6_io_vcsAvailable_0 )
  );
  VCRouterStateManagement VCRouterStateManagement_6(.clk(clk), .reset(reset),
       .io_inputBufferValid( RouterBuffer_6_io_deq_valid ),
       .io_routingComplete( R781 ),
       .io_inputBufferIsTail( T772 ),
       .io_vcAllocGranted( vcAllocator_io_resources_6_valid ),
       .io_swAllocGranted( T752 ),
       .io_creditsAvail( T733 ),
       .io_outputReady( T720 ),
       .io_currentState( VCRouterStateManagement_6_io_currentState )
  );
  ReplaceVCPort ReplaceVCPort_6(
       .io_oldFlit_x( T718 ),
       .io_newVCPort( T3133 ),
       .io_newFlit_x( ReplaceVCPort_6_io_newFlit_x )
  );
  Flit2FlitBundle Flit2FlitBundle_6(
       .io_inFlit_x( T712 )
       //.io_outHead_packetID(  )
       //.io_outHead_isTail(  )
       //.io_outHead_vcPort(  )
       //.io_outHead_packetType(  )
       //.io_outHead_destination_2(  )
       //.io_outHead_destination_1(  )
       //.io_outHead_destination_0(  )
       //.io_outHead_priorityLevel(  )
       //.io_outBody_packetID(  )
       //.io_outBody_isTail(  )
       //.io_outBody_vcPort(  )
       //.io_outBody_flitID(  )
       //.io_outBody_payload(  )
  );
  CreditGen CreditGen_7(
       .io_outCredit_grant( CreditGen_7_io_outCredit_grant ),
       .io_inGrant( T702 )
  );
  RouterRegFile RouterRegFile_7(.clk(clk), .reset(reset),
       .io_writeData( T700 ),
       .io_writeEnable( T697 ),
       //.io_full(  )
       .io_readData( RouterRegFile_7_io_readData ),
       .io_readValid( RouterRegFile_7_io_readValid ),
       .io_readIncrement( T684 ),
       .io_writePipelineReg_2( RouterRegFile_7_io_readPipelineReg_1 ),
       .io_writePipelineReg_1( RouterRegFile_7_io_readPipelineReg_0 ),
       .io_writePipelineReg_0( T3132 ),
       .io_wePipelineReg_2( T673 ),
       .io_wePipelineReg_1( T670 ),
       .io_wePipelineReg_0( T668 ),
       //.io_readPipelineReg_2(  )
       .io_readPipelineReg_1( RouterRegFile_7_io_readPipelineReg_1 ),
       .io_readPipelineReg_0( RouterRegFile_7_io_readPipelineReg_0 ),
       //.io_rvPipelineReg_2(  )
       .io_rvPipelineReg_1( RouterRegFile_7_io_rvPipelineReg_1 ),
       .io_rvPipelineReg_0( RouterRegFile_7_io_rvPipelineReg_0 )
  );
  RouterBuffer RouterBuffer_7(.clk(clk), .reset(reset),
       .io_enq_ready( RouterBuffer_7_io_enq_ready ),
       .io_enq_valid( T667 ),
       .io_enq_bits_x( io_inChannels_3_flit_x ),
       .io_deq_ready( T648 ),
       .io_deq_valid( RouterBuffer_7_io_deq_valid ),
       .io_deq_bits_x( RouterBuffer_7_io_deq_bits_x )
  );
  CMeshDOR_1 CMeshDOR_7(
       .io_inHeadFlit_packetID( T647 ),
       .io_inHeadFlit_isTail( T646 ),
       .io_inHeadFlit_vcPort( T645 ),
       .io_inHeadFlit_packetType( T644 ),
       .io_inHeadFlit_destination_2( T643 ),
       .io_inHeadFlit_destination_1( T642 ),
       .io_inHeadFlit_destination_0( T641 ),
       .io_inHeadFlit_priorityLevel( T638 ),
       .io_outHeadFlit_packetID( CMeshDOR_7_io_outHeadFlit_packetID ),
       .io_outHeadFlit_isTail( CMeshDOR_7_io_outHeadFlit_isTail ),
       .io_outHeadFlit_vcPort( CMeshDOR_7_io_outHeadFlit_vcPort ),
       .io_outHeadFlit_packetType( CMeshDOR_7_io_outHeadFlit_packetType ),
       .io_outHeadFlit_destination_2( CMeshDOR_7_io_outHeadFlit_destination_2 ),
       .io_outHeadFlit_destination_1( CMeshDOR_7_io_outHeadFlit_destination_1 ),
       .io_outHeadFlit_destination_0( CMeshDOR_7_io_outHeadFlit_destination_0 ),
       .io_outHeadFlit_priorityLevel( CMeshDOR_7_io_outHeadFlit_priorityLevel ),
       .io_result( CMeshDOR_7_io_result ),
       .io_vcsAvailable_4( CMeshDOR_7_io_vcsAvailable_4 ),
       .io_vcsAvailable_3( CMeshDOR_7_io_vcsAvailable_3 ),
       .io_vcsAvailable_2( CMeshDOR_7_io_vcsAvailable_2 ),
       .io_vcsAvailable_1( CMeshDOR_7_io_vcsAvailable_1 ),
       .io_vcsAvailable_0( CMeshDOR_7_io_vcsAvailable_0 )
  );
  VCRouterStateManagement VCRouterStateManagement_7(.clk(clk), .reset(reset),
       .io_inputBufferValid( RouterBuffer_7_io_deq_valid ),
       .io_routingComplete( R637 ),
       .io_inputBufferIsTail( T628 ),
       .io_vcAllocGranted( vcAllocator_io_resources_7_valid ),
       .io_swAllocGranted( T608 ),
       .io_creditsAvail( T589 ),
       .io_outputReady( T576 ),
       .io_currentState( VCRouterStateManagement_7_io_currentState )
  );
  ReplaceVCPort ReplaceVCPort_7(
       .io_oldFlit_x( T574 ),
       .io_newVCPort( T3126 ),
       .io_newFlit_x( ReplaceVCPort_7_io_newFlit_x )
  );
  Flit2FlitBundle Flit2FlitBundle_7(
       .io_inFlit_x( T568 )
       //.io_outHead_packetID(  )
       //.io_outHead_isTail(  )
       //.io_outHead_vcPort(  )
       //.io_outHead_packetType(  )
       //.io_outHead_destination_2(  )
       //.io_outHead_destination_1(  )
       //.io_outHead_destination_0(  )
       //.io_outHead_priorityLevel(  )
       //.io_outBody_packetID(  )
       //.io_outBody_isTail(  )
       //.io_outBody_vcPort(  )
       //.io_outBody_flitID(  )
       //.io_outBody_payload(  )
  );
  CreditGen CreditGen_8(
       .io_outCredit_grant( CreditGen_8_io_outCredit_grant ),
       .io_inGrant( T558 )
  );
  RouterRegFile RouterRegFile_8(.clk(clk), .reset(reset),
       .io_writeData( T556 ),
       .io_writeEnable( T553 ),
       //.io_full(  )
       .io_readData( RouterRegFile_8_io_readData ),
       .io_readValid( RouterRegFile_8_io_readValid ),
       .io_readIncrement( T540 ),
       .io_writePipelineReg_2( RouterRegFile_8_io_readPipelineReg_1 ),
       .io_writePipelineReg_1( RouterRegFile_8_io_readPipelineReg_0 ),
       .io_writePipelineReg_0( T3125 ),
       .io_wePipelineReg_2( T529 ),
       .io_wePipelineReg_1( T526 ),
       .io_wePipelineReg_0( T524 ),
       //.io_readPipelineReg_2(  )
       .io_readPipelineReg_1( RouterRegFile_8_io_readPipelineReg_1 ),
       .io_readPipelineReg_0( RouterRegFile_8_io_readPipelineReg_0 ),
       //.io_rvPipelineReg_2(  )
       .io_rvPipelineReg_1( RouterRegFile_8_io_rvPipelineReg_1 ),
       .io_rvPipelineReg_0( RouterRegFile_8_io_rvPipelineReg_0 )
  );
  RouterBuffer RouterBuffer_8(.clk(clk), .reset(reset),
       .io_enq_ready( RouterBuffer_8_io_enq_ready ),
       .io_enq_valid( T523 ),
       .io_enq_bits_x( io_inChannels_4_flit_x ),
       .io_deq_ready( T504 ),
       .io_deq_valid( RouterBuffer_8_io_deq_valid ),
       .io_deq_bits_x( RouterBuffer_8_io_deq_bits_x )
  );
  CMeshDOR_1 CMeshDOR_8(
       .io_inHeadFlit_packetID( T503 ),
       .io_inHeadFlit_isTail( T502 ),
       .io_inHeadFlit_vcPort( T501 ),
       .io_inHeadFlit_packetType( T500 ),
       .io_inHeadFlit_destination_2( T499 ),
       .io_inHeadFlit_destination_1( T498 ),
       .io_inHeadFlit_destination_0( T497 ),
       .io_inHeadFlit_priorityLevel( T494 ),
       .io_outHeadFlit_packetID( CMeshDOR_8_io_outHeadFlit_packetID ),
       .io_outHeadFlit_isTail( CMeshDOR_8_io_outHeadFlit_isTail ),
       .io_outHeadFlit_vcPort( CMeshDOR_8_io_outHeadFlit_vcPort ),
       .io_outHeadFlit_packetType( CMeshDOR_8_io_outHeadFlit_packetType ),
       .io_outHeadFlit_destination_2( CMeshDOR_8_io_outHeadFlit_destination_2 ),
       .io_outHeadFlit_destination_1( CMeshDOR_8_io_outHeadFlit_destination_1 ),
       .io_outHeadFlit_destination_0( CMeshDOR_8_io_outHeadFlit_destination_0 ),
       .io_outHeadFlit_priorityLevel( CMeshDOR_8_io_outHeadFlit_priorityLevel ),
       .io_result( CMeshDOR_8_io_result ),
       .io_vcsAvailable_4( CMeshDOR_8_io_vcsAvailable_4 ),
       .io_vcsAvailable_3( CMeshDOR_8_io_vcsAvailable_3 ),
       .io_vcsAvailable_2( CMeshDOR_8_io_vcsAvailable_2 ),
       .io_vcsAvailable_1( CMeshDOR_8_io_vcsAvailable_1 ),
       .io_vcsAvailable_0( CMeshDOR_8_io_vcsAvailable_0 )
  );
  VCRouterStateManagement VCRouterStateManagement_8(.clk(clk), .reset(reset),
       .io_inputBufferValid( RouterBuffer_8_io_deq_valid ),
       .io_routingComplete( R493 ),
       .io_inputBufferIsTail( T484 ),
       .io_vcAllocGranted( vcAllocator_io_resources_8_valid ),
       .io_swAllocGranted( T464 ),
       .io_creditsAvail( T445 ),
       .io_outputReady( T432 ),
       .io_currentState( VCRouterStateManagement_8_io_currentState )
  );
  ReplaceVCPort ReplaceVCPort_8(
       .io_oldFlit_x( T430 ),
       .io_newVCPort( T3119 ),
       .io_newFlit_x( ReplaceVCPort_8_io_newFlit_x )
  );
  Flit2FlitBundle Flit2FlitBundle_8(
       .io_inFlit_x( T424 )
       //.io_outHead_packetID(  )
       //.io_outHead_isTail(  )
       //.io_outHead_vcPort(  )
       //.io_outHead_packetType(  )
       //.io_outHead_destination_2(  )
       //.io_outHead_destination_1(  )
       //.io_outHead_destination_0(  )
       //.io_outHead_priorityLevel(  )
       //.io_outBody_packetID(  )
       //.io_outBody_isTail(  )
       //.io_outBody_vcPort(  )
       //.io_outBody_flitID(  )
       //.io_outBody_payload(  )
  );
  CreditGen CreditGen_9(
       .io_outCredit_grant( CreditGen_9_io_outCredit_grant ),
       .io_inGrant( T414 )
  );
  RouterRegFile RouterRegFile_9(.clk(clk), .reset(reset),
       .io_writeData( T412 ),
       .io_writeEnable( T409 ),
       //.io_full(  )
       .io_readData( RouterRegFile_9_io_readData ),
       .io_readValid( RouterRegFile_9_io_readValid ),
       .io_readIncrement( T396 ),
       .io_writePipelineReg_2( RouterRegFile_9_io_readPipelineReg_1 ),
       .io_writePipelineReg_1( RouterRegFile_9_io_readPipelineReg_0 ),
       .io_writePipelineReg_0( T3118 ),
       .io_wePipelineReg_2( T385 ),
       .io_wePipelineReg_1( T382 ),
       .io_wePipelineReg_0( T380 ),
       //.io_readPipelineReg_2(  )
       .io_readPipelineReg_1( RouterRegFile_9_io_readPipelineReg_1 ),
       .io_readPipelineReg_0( RouterRegFile_9_io_readPipelineReg_0 ),
       //.io_rvPipelineReg_2(  )
       .io_rvPipelineReg_1( RouterRegFile_9_io_rvPipelineReg_1 ),
       .io_rvPipelineReg_0( RouterRegFile_9_io_rvPipelineReg_0 )
  );
  RouterBuffer RouterBuffer_9(.clk(clk), .reset(reset),
       .io_enq_ready( RouterBuffer_9_io_enq_ready ),
       .io_enq_valid( T379 ),
       .io_enq_bits_x( io_inChannels_4_flit_x ),
       .io_deq_ready( T360 ),
       .io_deq_valid( RouterBuffer_9_io_deq_valid ),
       .io_deq_bits_x( RouterBuffer_9_io_deq_bits_x )
  );
  CMeshDOR_1 CMeshDOR_9(
       .io_inHeadFlit_packetID( T359 ),
       .io_inHeadFlit_isTail( T358 ),
       .io_inHeadFlit_vcPort( T357 ),
       .io_inHeadFlit_packetType( T356 ),
       .io_inHeadFlit_destination_2( T355 ),
       .io_inHeadFlit_destination_1( T354 ),
       .io_inHeadFlit_destination_0( T353 ),
       .io_inHeadFlit_priorityLevel( T350 ),
       .io_outHeadFlit_packetID( CMeshDOR_9_io_outHeadFlit_packetID ),
       .io_outHeadFlit_isTail( CMeshDOR_9_io_outHeadFlit_isTail ),
       .io_outHeadFlit_vcPort( CMeshDOR_9_io_outHeadFlit_vcPort ),
       .io_outHeadFlit_packetType( CMeshDOR_9_io_outHeadFlit_packetType ),
       .io_outHeadFlit_destination_2( CMeshDOR_9_io_outHeadFlit_destination_2 ),
       .io_outHeadFlit_destination_1( CMeshDOR_9_io_outHeadFlit_destination_1 ),
       .io_outHeadFlit_destination_0( CMeshDOR_9_io_outHeadFlit_destination_0 ),
       .io_outHeadFlit_priorityLevel( CMeshDOR_9_io_outHeadFlit_priorityLevel ),
       .io_result( CMeshDOR_9_io_result ),
       .io_vcsAvailable_4( CMeshDOR_9_io_vcsAvailable_4 ),
       .io_vcsAvailable_3( CMeshDOR_9_io_vcsAvailable_3 ),
       .io_vcsAvailable_2( CMeshDOR_9_io_vcsAvailable_2 ),
       .io_vcsAvailable_1( CMeshDOR_9_io_vcsAvailable_1 ),
       .io_vcsAvailable_0( CMeshDOR_9_io_vcsAvailable_0 )
  );
  VCRouterStateManagement VCRouterStateManagement_9(.clk(clk), .reset(reset),
       .io_inputBufferValid( RouterBuffer_9_io_deq_valid ),
       .io_routingComplete( R349 ),
       .io_inputBufferIsTail( T340 ),
       .io_vcAllocGranted( vcAllocator_io_resources_9_valid ),
       .io_swAllocGranted( T320 ),
       .io_creditsAvail( T301 ),
       .io_outputReady( T288 ),
       .io_currentState( VCRouterStateManagement_9_io_currentState )
  );
  ReplaceVCPort ReplaceVCPort_9(
       .io_oldFlit_x( T286 ),
       .io_newVCPort( T3112 ),
       .io_newFlit_x( ReplaceVCPort_9_io_newFlit_x )
  );
  Flit2FlitBundle Flit2FlitBundle_9(
       .io_inFlit_x( T280 )
       //.io_outHead_packetID(  )
       //.io_outHead_isTail(  )
       //.io_outHead_vcPort(  )
       //.io_outHead_packetType(  )
       //.io_outHead_destination_2(  )
       //.io_outHead_destination_1(  )
       //.io_outHead_destination_0(  )
       //.io_outHead_priorityLevel(  )
       //.io_outBody_packetID(  )
       //.io_outBody_isTail(  )
       //.io_outBody_vcPort(  )
       //.io_outBody_flitID(  )
       //.io_outBody_payload(  )
  );
  CreditCon CreditCon(.clk(clk), .reset(reset),
       .io_inCredit_grant( io_outChannels_0_credit_0_grant ),
       .io_inConsume( T278 ),
       .io_outCredit( CreditCon_io_outCredit )
       //.io_almostOut(  )
  );
  CreditCon CreditCon_1(.clk(clk), .reset(reset),
       .io_inCredit_grant( io_outChannels_0_credit_1_grant ),
       .io_inConsume( T268 ),
       .io_outCredit( CreditCon_1_io_outCredit )
       //.io_almostOut(  )
  );
  MuxN_1 MuxN(
       //.io_ins_1(  )
       //.io_ins_0(  )
       //.io_sel(  )
       //.io_out(  )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign MuxN.io_ins_1 = {1{1'b0}};
    assign MuxN.io_ins_0 = {1{1'b0}};
    assign MuxN.io_sel = {1{1'b0}};
// synthesis translate_on
`endif
  CreditCon CreditCon_2(.clk(clk), .reset(reset),
       .io_inCredit_grant( io_outChannels_1_credit_0_grant ),
       .io_inConsume( T266 ),
       .io_outCredit( CreditCon_2_io_outCredit )
       //.io_almostOut(  )
  );
  CreditCon CreditCon_3(.clk(clk), .reset(reset),
       .io_inCredit_grant( io_outChannels_1_credit_1_grant ),
       .io_inConsume( T256 ),
       .io_outCredit( CreditCon_3_io_outCredit )
       //.io_almostOut(  )
  );
  MuxN_1 MuxN_1(
       //.io_ins_1(  )
       //.io_ins_0(  )
       //.io_sel(  )
       //.io_out(  )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign MuxN_1.io_ins_1 = {1{1'b0}};
    assign MuxN_1.io_ins_0 = {1{1'b0}};
    assign MuxN_1.io_sel = {1{1'b0}};
// synthesis translate_on
`endif
  CreditCon CreditCon_4(.clk(clk), .reset(reset),
       .io_inCredit_grant( io_outChannels_2_credit_0_grant ),
       .io_inConsume( T254 ),
       .io_outCredit( CreditCon_4_io_outCredit )
       //.io_almostOut(  )
  );
  CreditCon CreditCon_5(.clk(clk), .reset(reset),
       .io_inCredit_grant( io_outChannels_2_credit_1_grant ),
       .io_inConsume( T244 ),
       .io_outCredit( CreditCon_5_io_outCredit )
       //.io_almostOut(  )
  );
  MuxN_1 MuxN_2(
       //.io_ins_1(  )
       //.io_ins_0(  )
       //.io_sel(  )
       //.io_out(  )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign MuxN_2.io_ins_1 = {1{1'b0}};
    assign MuxN_2.io_ins_0 = {1{1'b0}};
    assign MuxN_2.io_sel = {1{1'b0}};
// synthesis translate_on
`endif
  CreditCon CreditCon_6(.clk(clk), .reset(reset),
       .io_inCredit_grant( io_outChannels_3_credit_0_grant ),
       .io_inConsume( T242 ),
       .io_outCredit( CreditCon_6_io_outCredit )
       //.io_almostOut(  )
  );
  CreditCon CreditCon_7(.clk(clk), .reset(reset),
       .io_inCredit_grant( io_outChannels_3_credit_1_grant ),
       .io_inConsume( T232 ),
       .io_outCredit( CreditCon_7_io_outCredit )
       //.io_almostOut(  )
  );
  MuxN_1 MuxN_3(
       //.io_ins_1(  )
       //.io_ins_0(  )
       //.io_sel(  )
       //.io_out(  )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign MuxN_3.io_ins_1 = {1{1'b0}};
    assign MuxN_3.io_ins_0 = {1{1'b0}};
    assign MuxN_3.io_sel = {1{1'b0}};
// synthesis translate_on
`endif
  CreditCon CreditCon_8(.clk(clk), .reset(reset),
       .io_inCredit_grant( io_outChannels_4_credit_0_grant ),
       .io_inConsume( T230 ),
       .io_outCredit( CreditCon_8_io_outCredit )
       //.io_almostOut(  )
  );
  CreditCon CreditCon_9(.clk(clk), .reset(reset),
       .io_inCredit_grant( io_outChannels_4_credit_1_grant ),
       .io_inConsume( T220 ),
       .io_outCredit( CreditCon_9_io_outCredit )
       //.io_almostOut(  )
  );
  MuxN_1 MuxN_4(
       //.io_ins_1(  )
       //.io_ins_0(  )
       //.io_sel(  )
       //.io_out(  )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign MuxN_4.io_ins_1 = {1{1'b0}};
    assign MuxN_4.io_ins_0 = {1{1'b0}};
    assign MuxN_4.io_sel = {1{1'b0}};
// synthesis translate_on
`endif

  always @(posedge clk) begin
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T215 <= 1'b1;
  if(!T216 && T215 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "SimpleVCRouter: Flit with VC port/*? in < (class OpenSoC.SimpleVCRouter)>*/ Chisel.UInt(width=1, connect to 1 inputs: ([Chisel.Mux] in OpenSoC.SimpleVCRouter)) attempting to write to VC 0");
    $finish;
  end
// synthesis translate_on
`endif
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T198 <= 1'b1;
  if(!T199 && T198 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "SimpleVCRouter:Vector(1, 0) Insufficent space in input buffer - Credit Ready asserted when Routing In Buffer not ready inputPort= 0 curVC = 0");
    $finish;
  end
// synthesis translate_on
`endif
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T193 <= 1'b1;
  if(!T194 && T193 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "SimpleVCRouter: Flit with VC port/*? in < (class OpenSoC.SimpleVCRouter)>*/ Chisel.UInt(width=1, connect to 1 inputs: ([Chisel.Mux] in OpenSoC.SimpleVCRouter)) attempting to write to VC 1");
    $finish;
  end
// synthesis translate_on
`endif
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T176 <= 1'b1;
  if(!T177 && T176 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "SimpleVCRouter:Vector(1, 0) Insufficent space in input buffer - Credit Ready asserted when Routing In Buffer not ready inputPort= 0 curVC = 1");
    $finish;
  end
// synthesis translate_on
`endif
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T171 <= 1'b1;
  if(!T172 && T171 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "SimpleVCRouter: Flit with VC port/*? in < (class OpenSoC.SimpleVCRouter)>*/ Chisel.UInt(width=1, connect to 1 inputs: ([Chisel.Mux] in OpenSoC.SimpleVCRouter)) attempting to write to VC 0");
    $finish;
  end
// synthesis translate_on
`endif
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T154 <= 1'b1;
  if(!T155 && T154 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "SimpleVCRouter:Vector(1, 0) Insufficent space in input buffer - Credit Ready asserted when Routing In Buffer not ready inputPort= 1 curVC = 0");
    $finish;
  end
// synthesis translate_on
`endif
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T149 <= 1'b1;
  if(!T150 && T149 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "SimpleVCRouter: Flit with VC port/*? in < (class OpenSoC.SimpleVCRouter)>*/ Chisel.UInt(width=1, connect to 1 inputs: ([Chisel.Mux] in OpenSoC.SimpleVCRouter)) attempting to write to VC 1");
    $finish;
  end
// synthesis translate_on
`endif
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T132 <= 1'b1;
  if(!T133 && T132 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "SimpleVCRouter:Vector(1, 0) Insufficent space in input buffer - Credit Ready asserted when Routing In Buffer not ready inputPort= 1 curVC = 1");
    $finish;
  end
// synthesis translate_on
`endif
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T127 <= 1'b1;
  if(!T128 && T127 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "SimpleVCRouter: Flit with VC port/*? in < (class OpenSoC.SimpleVCRouter)>*/ Chisel.UInt(width=1, connect to 1 inputs: ([Chisel.Mux] in OpenSoC.SimpleVCRouter)) attempting to write to VC 0");
    $finish;
  end
// synthesis translate_on
`endif
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T110 <= 1'b1;
  if(!T111 && T110 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "SimpleVCRouter:Vector(1, 0) Insufficent space in input buffer - Credit Ready asserted when Routing In Buffer not ready inputPort= 2 curVC = 0");
    $finish;
  end
// synthesis translate_on
`endif
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T105 <= 1'b1;
  if(!T106 && T105 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "SimpleVCRouter: Flit with VC port/*? in < (class OpenSoC.SimpleVCRouter)>*/ Chisel.UInt(width=1, connect to 1 inputs: ([Chisel.Mux] in OpenSoC.SimpleVCRouter)) attempting to write to VC 1");
    $finish;
  end
// synthesis translate_on
`endif
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T88 <= 1'b1;
  if(!T89 && T88 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "SimpleVCRouter:Vector(1, 0) Insufficent space in input buffer - Credit Ready asserted when Routing In Buffer not ready inputPort= 2 curVC = 1");
    $finish;
  end
// synthesis translate_on
`endif
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T83 <= 1'b1;
  if(!T84 && T83 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "SimpleVCRouter: Flit with VC port/*? in < (class OpenSoC.SimpleVCRouter)>*/ Chisel.UInt(width=1, connect to 1 inputs: ([Chisel.Mux] in OpenSoC.SimpleVCRouter)) attempting to write to VC 0");
    $finish;
  end
// synthesis translate_on
`endif
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T66 <= 1'b1;
  if(!T67 && T66 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "SimpleVCRouter:Vector(1, 0) Insufficent space in input buffer - Credit Ready asserted when Routing In Buffer not ready inputPort= 3 curVC = 0");
    $finish;
  end
// synthesis translate_on
`endif
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T61 <= 1'b1;
  if(!T62 && T61 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "SimpleVCRouter: Flit with VC port/*? in < (class OpenSoC.SimpleVCRouter)>*/ Chisel.UInt(width=1, connect to 1 inputs: ([Chisel.Mux] in OpenSoC.SimpleVCRouter)) attempting to write to VC 1");
    $finish;
  end
// synthesis translate_on
`endif
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T44 <= 1'b1;
  if(!T45 && T44 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "SimpleVCRouter:Vector(1, 0) Insufficent space in input buffer - Credit Ready asserted when Routing In Buffer not ready inputPort= 3 curVC = 1");
    $finish;
  end
// synthesis translate_on
`endif
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T39 <= 1'b1;
  if(!T40 && T39 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "SimpleVCRouter: Flit with VC port/*? in < (class OpenSoC.SimpleVCRouter)>*/ Chisel.UInt(width=1, connect to 1 inputs: ([Chisel.Mux] in OpenSoC.SimpleVCRouter)) attempting to write to VC 0");
    $finish;
  end
// synthesis translate_on
`endif
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T22 <= 1'b1;
  if(!T23 && T22 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "SimpleVCRouter:Vector(1, 0) Insufficent space in input buffer - Credit Ready asserted when Routing In Buffer not ready inputPort= 4 curVC = 0");
    $finish;
  end
// synthesis translate_on
`endif
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T17 <= 1'b1;
  if(!T18 && T17 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "SimpleVCRouter: Flit with VC port/*? in < (class OpenSoC.SimpleVCRouter)>*/ Chisel.UInt(width=1, connect to 1 inputs: ([Chisel.Mux] in OpenSoC.SimpleVCRouter)) attempting to write to VC 1");
    $finish;
  end
// synthesis translate_on
`endif
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T0 <= 1'b1;
  if(!T1 && T0 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "SimpleVCRouter:Vector(1, 0) Insufficent space in input buffer - Credit Ready asserted when Routing In Buffer not ready inputPort= 4 curVC = 1");
    $finish;
  end
// synthesis translate_on
`endif
    if(reset) begin
      R282 <= 55'h0;
    end else if(T284) begin
      R282 <= T3114;
    end
    if(reset) begin
      R295 <= 3'h0;
    end else begin
      R295 <= CMeshDOR_9_io_result;
    end
    if(reset) begin
      R349 <= 1'h0;
    end else begin
      R349 <= RouterBuffer_9_io_deq_valid;
    end
    if(reset) begin
      R426 <= 55'h0;
    end else if(T428) begin
      R426 <= T3121;
    end
    if(reset) begin
      R439 <= 3'h0;
    end else begin
      R439 <= CMeshDOR_8_io_result;
    end
    if(reset) begin
      R493 <= 1'h0;
    end else begin
      R493 <= RouterBuffer_8_io_deq_valid;
    end
    if(reset) begin
      R570 <= 55'h0;
    end else if(T572) begin
      R570 <= T3128;
    end
    if(reset) begin
      R583 <= 3'h0;
    end else begin
      R583 <= CMeshDOR_7_io_result;
    end
    if(reset) begin
      R637 <= 1'h0;
    end else begin
      R637 <= RouterBuffer_7_io_deq_valid;
    end
    if(reset) begin
      R714 <= 55'h0;
    end else if(T716) begin
      R714 <= T3135;
    end
    if(reset) begin
      R727 <= 3'h0;
    end else begin
      R727 <= CMeshDOR_6_io_result;
    end
    if(reset) begin
      R781 <= 1'h0;
    end else begin
      R781 <= RouterBuffer_6_io_deq_valid;
    end
    if(reset) begin
      R858 <= 55'h0;
    end else if(T860) begin
      R858 <= T3142;
    end
    if(reset) begin
      R871 <= 3'h0;
    end else begin
      R871 <= CMeshDOR_5_io_result;
    end
    if(reset) begin
      R925 <= 1'h0;
    end else begin
      R925 <= RouterBuffer_5_io_deq_valid;
    end
    if(reset) begin
      R1002 <= 55'h0;
    end else if(T1004) begin
      R1002 <= T3149;
    end
    if(reset) begin
      R1015 <= 3'h0;
    end else begin
      R1015 <= CMeshDOR_4_io_result;
    end
    if(reset) begin
      R1069 <= 1'h0;
    end else begin
      R1069 <= RouterBuffer_4_io_deq_valid;
    end
    if(reset) begin
      R1146 <= 55'h0;
    end else if(T1148) begin
      R1146 <= T3156;
    end
    if(reset) begin
      R1159 <= 3'h0;
    end else begin
      R1159 <= CMeshDOR_3_io_result;
    end
    if(reset) begin
      R1213 <= 1'h0;
    end else begin
      R1213 <= RouterBuffer_3_io_deq_valid;
    end
    if(reset) begin
      R1290 <= 55'h0;
    end else if(T1292) begin
      R1290 <= T3163;
    end
    if(reset) begin
      R1303 <= 3'h0;
    end else begin
      R1303 <= CMeshDOR_2_io_result;
    end
    if(reset) begin
      R1357 <= 1'h0;
    end else begin
      R1357 <= RouterBuffer_2_io_deq_valid;
    end
    if(reset) begin
      R1434 <= 55'h0;
    end else if(T1436) begin
      R1434 <= T3170;
    end
    if(reset) begin
      R1447 <= 3'h0;
    end else begin
      R1447 <= CMeshDOR_1_io_result;
    end
    if(reset) begin
      R1501 <= 1'h0;
    end else begin
      R1501 <= RouterBuffer_1_io_deq_valid;
    end
    if(reset) begin
      R1578 <= 55'h0;
    end else if(T1580) begin
      R1578 <= T3177;
    end
    if(reset) begin
      R1591 <= 3'h0;
    end else begin
      R1591 <= CMeshDOR_io_result;
    end
    if(reset) begin
      R1645 <= 1'h0;
    end else begin
      R1645 <= RouterBuffer_io_deq_valid;
    end
    validVCs_0_0 <= CMeshDOR_io_vcsAvailable_0;
    R2176 <= T2177;
    R2181 <= T2182;
    validVCs_0_1 <= CMeshDOR_io_vcsAvailable_1;
    R2186 <= T2187;
    R2191 <= T2192;
    validVCs_0_2 <= CMeshDOR_io_vcsAvailable_2;
    R2196 <= T2197;
    R2201 <= T2202;
    validVCs_0_3 <= CMeshDOR_io_vcsAvailable_3;
    R2206 <= T2207;
    R2211 <= T2212;
    validVCs_0_4 <= CMeshDOR_io_vcsAvailable_4;
    R2216 <= T2217;
    R2221 <= T2222;
    validVCs_1_0 <= CMeshDOR_1_io_vcsAvailable_0;
    R2226 <= T2227;
    R2231 <= T2232;
    validVCs_1_1 <= CMeshDOR_1_io_vcsAvailable_1;
    R2236 <= T2237;
    R2241 <= T2242;
    validVCs_1_2 <= CMeshDOR_1_io_vcsAvailable_2;
    R2246 <= T2247;
    R2251 <= T2252;
    validVCs_1_3 <= CMeshDOR_1_io_vcsAvailable_3;
    R2256 <= T2257;
    R2261 <= T2262;
    validVCs_1_4 <= CMeshDOR_1_io_vcsAvailable_4;
    R2266 <= T2267;
    R2271 <= T2272;
    validVCs_2_0 <= CMeshDOR_2_io_vcsAvailable_0;
    R2276 <= T2277;
    R2281 <= T2282;
    validVCs_2_1 <= CMeshDOR_2_io_vcsAvailable_1;
    R2286 <= T2287;
    R2291 <= T2292;
    validVCs_2_2 <= CMeshDOR_2_io_vcsAvailable_2;
    R2296 <= T2297;
    R2301 <= T2302;
    validVCs_2_3 <= CMeshDOR_2_io_vcsAvailable_3;
    R2306 <= T2307;
    R2311 <= T2312;
    validVCs_2_4 <= CMeshDOR_2_io_vcsAvailable_4;
    R2316 <= T2317;
    R2321 <= T2322;
    validVCs_3_0 <= CMeshDOR_3_io_vcsAvailable_0;
    R2326 <= T2327;
    R2331 <= T2332;
    validVCs_3_1 <= CMeshDOR_3_io_vcsAvailable_1;
    R2336 <= T2337;
    R2341 <= T2342;
    validVCs_3_2 <= CMeshDOR_3_io_vcsAvailable_2;
    R2346 <= T2347;
    R2351 <= T2352;
    validVCs_3_3 <= CMeshDOR_3_io_vcsAvailable_3;
    R2356 <= T2357;
    R2361 <= T2362;
    validVCs_3_4 <= CMeshDOR_3_io_vcsAvailable_4;
    R2366 <= T2367;
    R2371 <= T2372;
    validVCs_4_0 <= CMeshDOR_4_io_vcsAvailable_0;
    R2376 <= T2377;
    R2381 <= T2382;
    validVCs_4_1 <= CMeshDOR_4_io_vcsAvailable_1;
    R2386 <= T2387;
    R2391 <= T2392;
    validVCs_4_2 <= CMeshDOR_4_io_vcsAvailable_2;
    R2396 <= T2397;
    R2401 <= T2402;
    validVCs_4_3 <= CMeshDOR_4_io_vcsAvailable_3;
    R2406 <= T2407;
    R2411 <= T2412;
    validVCs_4_4 <= CMeshDOR_4_io_vcsAvailable_4;
    R2416 <= T2417;
    R2421 <= T2422;
    validVCs_5_0 <= CMeshDOR_5_io_vcsAvailable_0;
    R2426 <= T2427;
    R2431 <= T2432;
    validVCs_5_1 <= CMeshDOR_5_io_vcsAvailable_1;
    R2436 <= T2437;
    R2441 <= T2442;
    validVCs_5_2 <= CMeshDOR_5_io_vcsAvailable_2;
    R2446 <= T2447;
    R2451 <= T2452;
    validVCs_5_3 <= CMeshDOR_5_io_vcsAvailable_3;
    R2456 <= T2457;
    R2461 <= T2462;
    validVCs_5_4 <= CMeshDOR_5_io_vcsAvailable_4;
    R2466 <= T2467;
    R2471 <= T2472;
    validVCs_6_0 <= CMeshDOR_6_io_vcsAvailable_0;
    R2476 <= T2477;
    R2481 <= T2482;
    validVCs_6_1 <= CMeshDOR_6_io_vcsAvailable_1;
    R2486 <= T2487;
    R2491 <= T2492;
    validVCs_6_2 <= CMeshDOR_6_io_vcsAvailable_2;
    R2496 <= T2497;
    R2501 <= T2502;
    validVCs_6_3 <= CMeshDOR_6_io_vcsAvailable_3;
    R2506 <= T2507;
    R2511 <= T2512;
    validVCs_6_4 <= CMeshDOR_6_io_vcsAvailable_4;
    R2516 <= T2517;
    R2521 <= T2522;
    validVCs_7_0 <= CMeshDOR_7_io_vcsAvailable_0;
    R2526 <= T2527;
    R2531 <= T2532;
    validVCs_7_1 <= CMeshDOR_7_io_vcsAvailable_1;
    R2536 <= T2537;
    R2541 <= T2542;
    validVCs_7_2 <= CMeshDOR_7_io_vcsAvailable_2;
    R2546 <= T2547;
    R2551 <= T2552;
    validVCs_7_3 <= CMeshDOR_7_io_vcsAvailable_3;
    R2556 <= T2557;
    R2561 <= T2562;
    validVCs_7_4 <= CMeshDOR_7_io_vcsAvailable_4;
    R2566 <= T2567;
    R2571 <= T2572;
    validVCs_8_0 <= CMeshDOR_8_io_vcsAvailable_0;
    R2576 <= T2577;
    R2581 <= T2582;
    validVCs_8_1 <= CMeshDOR_8_io_vcsAvailable_1;
    R2586 <= T2587;
    R2591 <= T2592;
    validVCs_8_2 <= CMeshDOR_8_io_vcsAvailable_2;
    R2596 <= T2597;
    R2601 <= T2602;
    validVCs_8_3 <= CMeshDOR_8_io_vcsAvailable_3;
    R2606 <= T2607;
    R2611 <= T2612;
    validVCs_8_4 <= CMeshDOR_8_io_vcsAvailable_4;
    R2616 <= T2617;
    R2621 <= T2622;
    validVCs_9_0 <= CMeshDOR_9_io_vcsAvailable_0;
    R2626 <= T2627;
    R2631 <= T2632;
    validVCs_9_1 <= CMeshDOR_9_io_vcsAvailable_1;
    R2636 <= T2637;
    R2641 <= T2642;
    validVCs_9_2 <= CMeshDOR_9_io_vcsAvailable_2;
    R2646 <= T2647;
    R2651 <= T2652;
    validVCs_9_3 <= CMeshDOR_9_io_vcsAvailable_3;
    R2656 <= T2657;
    R2661 <= T2662;
    validVCs_9_4 <= CMeshDOR_9_io_vcsAvailable_4;
    R2666 <= T2667;
    R2671 <= T2672;
    if(reset) begin
      R2675 <= 3'h0;
    end else if(T1670) begin
      R2675 <= T2677;
    end
    if(reset) begin
      R2683 <= 8'h0;
    end else begin
      R2683 <= T2684;
    end
    if(reset) begin
      R2688 <= 1'h1;
    end else begin
      R2688 <= T1692;
    end
    if(reset) begin
      R2689 <= 3'h0;
    end else if(T1526) begin
      R2689 <= T2691;
    end
    if(reset) begin
      R2697 <= 8'h0;
    end else begin
      R2697 <= T2698;
    end
    if(reset) begin
      R2702 <= 1'h1;
    end else begin
      R2702 <= T1548;
    end
    if(reset) begin
      R2703 <= 3'h0;
    end else if(T1382) begin
      R2703 <= T2705;
    end
    if(reset) begin
      R2711 <= 8'h0;
    end else begin
      R2711 <= T2712;
    end
    if(reset) begin
      R2716 <= 1'h1;
    end else begin
      R2716 <= T1404;
    end
    if(reset) begin
      R2717 <= 3'h0;
    end else if(T1238) begin
      R2717 <= T2719;
    end
    if(reset) begin
      R2725 <= 8'h0;
    end else begin
      R2725 <= T2726;
    end
    if(reset) begin
      R2730 <= 1'h1;
    end else begin
      R2730 <= T1260;
    end
    if(reset) begin
      R2731 <= 3'h0;
    end else if(T1094) begin
      R2731 <= T2733;
    end
    if(reset) begin
      R2739 <= 8'h0;
    end else begin
      R2739 <= T2740;
    end
    if(reset) begin
      R2744 <= 1'h1;
    end else begin
      R2744 <= T1116;
    end
    if(reset) begin
      R2745 <= 3'h0;
    end else if(T950) begin
      R2745 <= T2747;
    end
    if(reset) begin
      R2753 <= 8'h0;
    end else begin
      R2753 <= T2754;
    end
    if(reset) begin
      R2758 <= 1'h1;
    end else begin
      R2758 <= T972;
    end
    if(reset) begin
      R2759 <= 3'h0;
    end else if(T806) begin
      R2759 <= T2761;
    end
    if(reset) begin
      R2767 <= 8'h0;
    end else begin
      R2767 <= T2768;
    end
    if(reset) begin
      R2772 <= 1'h1;
    end else begin
      R2772 <= T828;
    end
    if(reset) begin
      R2773 <= 3'h0;
    end else if(T662) begin
      R2773 <= T2775;
    end
    if(reset) begin
      R2781 <= 8'h0;
    end else begin
      R2781 <= T2782;
    end
    if(reset) begin
      R2786 <= 1'h1;
    end else begin
      R2786 <= T684;
    end
    if(reset) begin
      R2787 <= 3'h0;
    end else if(T518) begin
      R2787 <= T2789;
    end
    if(reset) begin
      R2795 <= 8'h0;
    end else begin
      R2795 <= T2796;
    end
    if(reset) begin
      R2800 <= 1'h1;
    end else begin
      R2800 <= T540;
    end
    if(reset) begin
      R2801 <= 3'h0;
    end else if(T374) begin
      R2801 <= T2803;
    end
    if(reset) begin
      R2809 <= 8'h0;
    end else begin
      R2809 <= T2810;
    end
    if(reset) begin
      R2814 <= 1'h1;
    end else begin
      R2814 <= T396;
    end
    R3097 <= T2094;
    if(reset) begin
      R3098 <= T3099;
    end else begin
      R3098 <= switch_io_outPorts_0_x;
    end
    R3100 <= T2031;
    if(reset) begin
      R3101 <= T3102;
    end else begin
      R3101 <= switch_io_outPorts_1_x;
    end
    R3103 <= T1968;
    if(reset) begin
      R3104 <= T3105;
    end else begin
      R3104 <= switch_io_outPorts_2_x;
    end
    R3106 <= T1905;
    if(reset) begin
      R3107 <= T3108;
    end else begin
      R3107 <= switch_io_outPorts_3_x;
    end
    R3109 <= T1722;
    if(reset) begin
      R3110 <= T3111;
    end else begin
      R3110 <= switch_io_outPorts_4_x;
    end
  end
endmodule

module VCRouterWrapper_1(input clk, input reset,
    input [54:0] io_inChannels_4_flit_x,
    input  io_inChannels_4_flitValid,
    output io_inChannels_4_credit_1_grant,
    output io_inChannels_4_credit_0_grant,
    input [54:0] io_inChannels_3_flit_x,
    input  io_inChannels_3_flitValid,
    output io_inChannels_3_credit_1_grant,
    output io_inChannels_3_credit_0_grant,
    input [54:0] io_inChannels_2_flit_x,
    input  io_inChannels_2_flitValid,
    output io_inChannels_2_credit_1_grant,
    output io_inChannels_2_credit_0_grant,
    input [54:0] io_inChannels_1_flit_x,
    input  io_inChannels_1_flitValid,
    output io_inChannels_1_credit_1_grant,
    output io_inChannels_1_credit_0_grant,
    input [54:0] io_inChannels_0_flit_x,
    input  io_inChannels_0_flitValid,
    output io_inChannels_0_credit_1_grant,
    output io_inChannels_0_credit_0_grant,
    output[54:0] io_outChannels_4_flit_x,
    output io_outChannels_4_flitValid,
    input  io_outChannels_4_credit_1_grant,
    input  io_outChannels_4_credit_0_grant,
    output[54:0] io_outChannels_3_flit_x,
    output io_outChannels_3_flitValid,
    input  io_outChannels_3_credit_1_grant,
    input  io_outChannels_3_credit_0_grant,
    output[54:0] io_outChannels_2_flit_x,
    output io_outChannels_2_flitValid,
    input  io_outChannels_2_credit_1_grant,
    input  io_outChannels_2_credit_0_grant,
    output[54:0] io_outChannels_1_flit_x,
    output io_outChannels_1_flitValid,
    input  io_outChannels_1_credit_1_grant,
    input  io_outChannels_1_credit_0_grant,
    output[54:0] io_outChannels_0_flit_x,
    output io_outChannels_0_flitValid,
    input  io_outChannels_0_credit_1_grant,
    input  io_outChannels_0_credit_0_grant,
    output[31:0] io_counters_1_counterVal,
    output[7:0] io_counters_1_counterIndex,
    output[31:0] io_counters_0_counterVal,
    output[7:0] io_counters_0_counterIndex,
    input  io_bypass
);

  wire bp_io_x_inChannels_4_credit_1_grant;
  wire bp_io_x_inChannels_4_credit_0_grant;
  wire bp_io_x_inChannels_3_credit_1_grant;
  wire bp_io_x_inChannels_3_credit_0_grant;
  wire bp_io_x_inChannels_2_credit_1_grant;
  wire bp_io_x_inChannels_2_credit_0_grant;
  wire bp_io_x_inChannels_1_credit_1_grant;
  wire bp_io_x_inChannels_1_credit_0_grant;
  wire bp_io_x_inChannels_0_credit_1_grant;
  wire bp_io_x_inChannels_0_credit_0_grant;
  wire[54:0] bp_io_x_outChannels_4_flit_x;
  wire bp_io_x_outChannels_4_flitValid;
  wire[54:0] bp_io_x_outChannels_3_flit_x;
  wire bp_io_x_outChannels_3_flitValid;
  wire[54:0] bp_io_x_outChannels_2_flit_x;
  wire bp_io_x_outChannels_2_flitValid;
  wire[54:0] bp_io_x_outChannels_1_flit_x;
  wire bp_io_x_outChannels_1_flitValid;
  wire[54:0] bp_io_x_outChannels_0_flit_x;
  wire bp_io_x_outChannels_0_flitValid;
  wire[31:0] bp_io_x_counters_1_counterVal;
  wire[7:0] bp_io_x_counters_1_counterIndex;
  wire[31:0] bp_io_x_counters_0_counterVal;
  wire[7:0] bp_io_x_counters_0_counterIndex;
  wire[54:0] bp_io_y_inChannels_4_flit_x;
  wire bp_io_y_inChannels_4_flitValid;
  wire[54:0] bp_io_y_inChannels_3_flit_x;
  wire bp_io_y_inChannels_3_flitValid;
  wire[54:0] bp_io_y_inChannels_2_flit_x;
  wire bp_io_y_inChannels_2_flitValid;
  wire[54:0] bp_io_y_inChannels_1_flit_x;
  wire bp_io_y_inChannels_1_flitValid;
  wire[54:0] bp_io_y_inChannels_0_flit_x;
  wire bp_io_y_inChannels_0_flitValid;
  wire bp_io_y_outChannels_4_credit_1_grant;
  wire bp_io_y_outChannels_4_credit_0_grant;
  wire bp_io_y_outChannels_3_credit_1_grant;
  wire bp_io_y_outChannels_3_credit_0_grant;
  wire bp_io_y_outChannels_2_credit_1_grant;
  wire bp_io_y_outChannels_2_credit_0_grant;
  wire bp_io_y_outChannels_1_credit_1_grant;
  wire bp_io_y_outChannels_1_credit_0_grant;
  wire bp_io_y_outChannels_0_credit_1_grant;
  wire bp_io_y_outChannels_0_credit_0_grant;
  wire x_io_inChannels_4_credit_1_grant;
  wire x_io_inChannels_4_credit_0_grant;
  wire x_io_inChannels_3_credit_1_grant;
  wire x_io_inChannels_3_credit_0_grant;
  wire x_io_inChannels_2_credit_1_grant;
  wire x_io_inChannels_2_credit_0_grant;
  wire x_io_inChannels_1_credit_1_grant;
  wire x_io_inChannels_1_credit_0_grant;
  wire x_io_inChannels_0_credit_1_grant;
  wire x_io_inChannels_0_credit_0_grant;
  wire[54:0] x_io_outChannels_4_flit_x;
  wire x_io_outChannels_4_flitValid;
  wire[54:0] x_io_outChannels_3_flit_x;
  wire x_io_outChannels_3_flitValid;
  wire[54:0] x_io_outChannels_2_flit_x;
  wire x_io_outChannels_2_flitValid;
  wire[54:0] x_io_outChannels_1_flit_x;
  wire x_io_outChannels_1_flitValid;
  wire[54:0] x_io_outChannels_0_flit_x;
  wire x_io_outChannels_0_flitValid;
  wire[31:0] x_io_counters_0_counterVal;


  assign io_counters_0_counterIndex = bp_io_x_counters_0_counterIndex;
  assign io_counters_0_counterVal = bp_io_x_counters_0_counterVal;
  assign io_counters_1_counterIndex = bp_io_x_counters_1_counterIndex;
  assign io_counters_1_counterVal = bp_io_x_counters_1_counterVal;
  assign io_outChannels_0_flitValid = bp_io_x_outChannels_0_flitValid;
  assign io_outChannels_0_flit_x = bp_io_x_outChannels_0_flit_x;
  assign io_outChannels_1_flitValid = bp_io_x_outChannels_1_flitValid;
  assign io_outChannels_1_flit_x = bp_io_x_outChannels_1_flit_x;
  assign io_outChannels_2_flitValid = bp_io_x_outChannels_2_flitValid;
  assign io_outChannels_2_flit_x = bp_io_x_outChannels_2_flit_x;
  assign io_outChannels_3_flitValid = bp_io_x_outChannels_3_flitValid;
  assign io_outChannels_3_flit_x = bp_io_x_outChannels_3_flit_x;
  assign io_outChannels_4_flitValid = bp_io_x_outChannels_4_flitValid;
  assign io_outChannels_4_flit_x = bp_io_x_outChannels_4_flit_x;
  assign io_inChannels_0_credit_0_grant = bp_io_x_inChannels_0_credit_0_grant;
  assign io_inChannels_0_credit_1_grant = bp_io_x_inChannels_0_credit_1_grant;
  assign io_inChannels_1_credit_0_grant = bp_io_x_inChannels_1_credit_0_grant;
  assign io_inChannels_1_credit_1_grant = bp_io_x_inChannels_1_credit_1_grant;
  assign io_inChannels_2_credit_0_grant = bp_io_x_inChannels_2_credit_0_grant;
  assign io_inChannels_2_credit_1_grant = bp_io_x_inChannels_2_credit_1_grant;
  assign io_inChannels_3_credit_0_grant = bp_io_x_inChannels_3_credit_0_grant;
  assign io_inChannels_3_credit_1_grant = bp_io_x_inChannels_3_credit_1_grant;
  assign io_inChannels_4_credit_0_grant = bp_io_x_inChannels_4_credit_0_grant;
  assign io_inChannels_4_credit_1_grant = bp_io_x_inChannels_4_credit_1_grant;
  wire clkOut;
  VCRouterBypass bp(.clk(clk), .reset(reset),
       .io_x_inChannels_4_flit_x( io_inChannels_4_flit_x ),
       .io_x_inChannels_4_flitValid( io_inChannels_4_flitValid ),
       .io_x_inChannels_4_credit_1_grant( bp_io_x_inChannels_4_credit_1_grant ),
       .io_x_inChannels_4_credit_0_grant( bp_io_x_inChannels_4_credit_0_grant ),
       .io_x_inChannels_3_flit_x( io_inChannels_3_flit_x ),
       .io_x_inChannels_3_flitValid( io_inChannels_3_flitValid ),
       .io_x_inChannels_3_credit_1_grant( bp_io_x_inChannels_3_credit_1_grant ),
       .io_x_inChannels_3_credit_0_grant( bp_io_x_inChannels_3_credit_0_grant ),
       .io_x_inChannels_2_flit_x( io_inChannels_2_flit_x ),
       .io_x_inChannels_2_flitValid( io_inChannels_2_flitValid ),
       .io_x_inChannels_2_credit_1_grant( bp_io_x_inChannels_2_credit_1_grant ),
       .io_x_inChannels_2_credit_0_grant( bp_io_x_inChannels_2_credit_0_grant ),
       .io_x_inChannels_1_flit_x( io_inChannels_1_flit_x ),
       .io_x_inChannels_1_flitValid( io_inChannels_1_flitValid ),
       .io_x_inChannels_1_credit_1_grant( bp_io_x_inChannels_1_credit_1_grant ),
       .io_x_inChannels_1_credit_0_grant( bp_io_x_inChannels_1_credit_0_grant ),
       .io_x_inChannels_0_flit_x( io_inChannels_0_flit_x ),
       .io_x_inChannels_0_flitValid( io_inChannels_0_flitValid ),
       .io_x_inChannels_0_credit_1_grant( bp_io_x_inChannels_0_credit_1_grant ),
       .io_x_inChannels_0_credit_0_grant( bp_io_x_inChannels_0_credit_0_grant ),
       .io_x_outChannels_4_flit_x( bp_io_x_outChannels_4_flit_x ),
       .io_x_outChannels_4_flitValid( bp_io_x_outChannels_4_flitValid ),
       .io_x_outChannels_4_credit_1_grant( io_outChannels_4_credit_1_grant ),
       .io_x_outChannels_4_credit_0_grant( io_outChannels_4_credit_0_grant ),
       .io_x_outChannels_3_flit_x( bp_io_x_outChannels_3_flit_x ),
       .io_x_outChannels_3_flitValid( bp_io_x_outChannels_3_flitValid ),
       .io_x_outChannels_3_credit_1_grant( io_outChannels_3_credit_1_grant ),
       .io_x_outChannels_3_credit_0_grant( io_outChannels_3_credit_0_grant ),
       .io_x_outChannels_2_flit_x( bp_io_x_outChannels_2_flit_x ),
       .io_x_outChannels_2_flitValid( bp_io_x_outChannels_2_flitValid ),
       .io_x_outChannels_2_credit_1_grant( io_outChannels_2_credit_1_grant ),
       .io_x_outChannels_2_credit_0_grant( io_outChannels_2_credit_0_grant ),
       .io_x_outChannels_1_flit_x( bp_io_x_outChannels_1_flit_x ),
       .io_x_outChannels_1_flitValid( bp_io_x_outChannels_1_flitValid ),
       .io_x_outChannels_1_credit_1_grant( io_outChannels_1_credit_1_grant ),
       .io_x_outChannels_1_credit_0_grant( io_outChannels_1_credit_0_grant ),
       .io_x_outChannels_0_flit_x( bp_io_x_outChannels_0_flit_x ),
       .io_x_outChannels_0_flitValid( bp_io_x_outChannels_0_flitValid ),
       .io_x_outChannels_0_credit_1_grant( io_outChannels_0_credit_1_grant ),
       .io_x_outChannels_0_credit_0_grant( io_outChannels_0_credit_0_grant ),
       .io_x_counters_1_counterVal( bp_io_x_counters_1_counterVal ),
       .io_x_counters_1_counterIndex( bp_io_x_counters_1_counterIndex ),
       .io_x_counters_0_counterVal( bp_io_x_counters_0_counterVal ),
       .io_x_counters_0_counterIndex( bp_io_x_counters_0_counterIndex ),
       .io_y_inChannels_4_flit_x( bp_io_y_inChannels_4_flit_x ),
       .io_y_inChannels_4_flitValid( bp_io_y_inChannels_4_flitValid ),
       .io_y_inChannels_4_credit_1_grant( x_io_inChannels_4_credit_1_grant ),
       .io_y_inChannels_4_credit_0_grant( x_io_inChannels_4_credit_0_grant ),
       .io_y_inChannels_3_flit_x( bp_io_y_inChannels_3_flit_x ),
       .io_y_inChannels_3_flitValid( bp_io_y_inChannels_3_flitValid ),
       .io_y_inChannels_3_credit_1_grant( x_io_inChannels_3_credit_1_grant ),
       .io_y_inChannels_3_credit_0_grant( x_io_inChannels_3_credit_0_grant ),
       .io_y_inChannels_2_flit_x( bp_io_y_inChannels_2_flit_x ),
       .io_y_inChannels_2_flitValid( bp_io_y_inChannels_2_flitValid ),
       .io_y_inChannels_2_credit_1_grant( x_io_inChannels_2_credit_1_grant ),
       .io_y_inChannels_2_credit_0_grant( x_io_inChannels_2_credit_0_grant ),
       .io_y_inChannels_1_flit_x( bp_io_y_inChannels_1_flit_x ),
       .io_y_inChannels_1_flitValid( bp_io_y_inChannels_1_flitValid ),
       .io_y_inChannels_1_credit_1_grant( x_io_inChannels_1_credit_1_grant ),
       .io_y_inChannels_1_credit_0_grant( x_io_inChannels_1_credit_0_grant ),
       .io_y_inChannels_0_flit_x( bp_io_y_inChannels_0_flit_x ),
       .io_y_inChannels_0_flitValid( bp_io_y_inChannels_0_flitValid ),
       .io_y_inChannels_0_credit_1_grant( x_io_inChannels_0_credit_1_grant ),
       .io_y_inChannels_0_credit_0_grant( x_io_inChannels_0_credit_0_grant ),
       .io_y_outChannels_4_flit_x( x_io_outChannels_4_flit_x ),
       .io_y_outChannels_4_flitValid( x_io_outChannels_4_flitValid ),
       .io_y_outChannels_4_credit_1_grant( bp_io_y_outChannels_4_credit_1_grant ),
       .io_y_outChannels_4_credit_0_grant( bp_io_y_outChannels_4_credit_0_grant ),
       .io_y_outChannels_3_flit_x( x_io_outChannels_3_flit_x ),
       .io_y_outChannels_3_flitValid( x_io_outChannels_3_flitValid ),
       .io_y_outChannels_3_credit_1_grant( bp_io_y_outChannels_3_credit_1_grant ),
       .io_y_outChannels_3_credit_0_grant( bp_io_y_outChannels_3_credit_0_grant ),
       .io_y_outChannels_2_flit_x( x_io_outChannels_2_flit_x ),
       .io_y_outChannels_2_flitValid( x_io_outChannels_2_flitValid ),
       .io_y_outChannels_2_credit_1_grant( bp_io_y_outChannels_2_credit_1_grant ),
       .io_y_outChannels_2_credit_0_grant( bp_io_y_outChannels_2_credit_0_grant ),
       .io_y_outChannels_1_flit_x( x_io_outChannels_1_flit_x ),
       .io_y_outChannels_1_flitValid( x_io_outChannels_1_flitValid ),
       .io_y_outChannels_1_credit_1_grant( bp_io_y_outChannels_1_credit_1_grant ),
       .io_y_outChannels_1_credit_0_grant( bp_io_y_outChannels_1_credit_0_grant ),
       .io_y_outChannels_0_flit_x( x_io_outChannels_0_flit_x ),
       .io_y_outChannels_0_flitValid( x_io_outChannels_0_flitValid ),
       .io_y_outChannels_0_credit_1_grant( bp_io_y_outChannels_0_credit_1_grant ),
       .io_y_outChannels_0_credit_0_grant( bp_io_y_outChannels_0_credit_0_grant ),
       //.io_y_counters_1_counterVal(  )
       //.io_y_counters_1_counterIndex(  )
       .io_y_counters_0_counterVal( x_io_counters_0_counterVal ),
       //.io_y_counters_0_counterIndex(  )
       .io_bypass( io_bypass ),
       .io_clkOut(clkOut)
  );
  SimpleVCRouter_1 x(.clk(clkOut), .reset(reset),
       .io_inChannels_4_flit_x( bp_io_y_inChannels_4_flit_x ),
       .io_inChannels_4_flitValid( bp_io_y_inChannels_4_flitValid ),
       .io_inChannels_4_credit_1_grant( x_io_inChannels_4_credit_1_grant ),
       .io_inChannels_4_credit_0_grant( x_io_inChannels_4_credit_0_grant ),
       .io_inChannels_3_flit_x( bp_io_y_inChannels_3_flit_x ),
       .io_inChannels_3_flitValid( bp_io_y_inChannels_3_flitValid ),
       .io_inChannels_3_credit_1_grant( x_io_inChannels_3_credit_1_grant ),
       .io_inChannels_3_credit_0_grant( x_io_inChannels_3_credit_0_grant ),
       .io_inChannels_2_flit_x( bp_io_y_inChannels_2_flit_x ),
       .io_inChannels_2_flitValid( bp_io_y_inChannels_2_flitValid ),
       .io_inChannels_2_credit_1_grant( x_io_inChannels_2_credit_1_grant ),
       .io_inChannels_2_credit_0_grant( x_io_inChannels_2_credit_0_grant ),
       .io_inChannels_1_flit_x( bp_io_y_inChannels_1_flit_x ),
       .io_inChannels_1_flitValid( bp_io_y_inChannels_1_flitValid ),
       .io_inChannels_1_credit_1_grant( x_io_inChannels_1_credit_1_grant ),
       .io_inChannels_1_credit_0_grant( x_io_inChannels_1_credit_0_grant ),
       .io_inChannels_0_flit_x( bp_io_y_inChannels_0_flit_x ),
       .io_inChannels_0_flitValid( bp_io_y_inChannels_0_flitValid ),
       .io_inChannels_0_credit_1_grant( x_io_inChannels_0_credit_1_grant ),
       .io_inChannels_0_credit_0_grant( x_io_inChannels_0_credit_0_grant ),
       .io_outChannels_4_flit_x( x_io_outChannels_4_flit_x ),
       .io_outChannels_4_flitValid( x_io_outChannels_4_flitValid ),
       .io_outChannels_4_credit_1_grant( bp_io_y_outChannels_4_credit_1_grant ),
       .io_outChannels_4_credit_0_grant( bp_io_y_outChannels_4_credit_0_grant ),
       .io_outChannels_3_flit_x( x_io_outChannels_3_flit_x ),
       .io_outChannels_3_flitValid( x_io_outChannels_3_flitValid ),
       .io_outChannels_3_credit_1_grant( bp_io_y_outChannels_3_credit_1_grant ),
       .io_outChannels_3_credit_0_grant( bp_io_y_outChannels_3_credit_0_grant ),
       .io_outChannels_2_flit_x( x_io_outChannels_2_flit_x ),
       .io_outChannels_2_flitValid( x_io_outChannels_2_flitValid ),
       .io_outChannels_2_credit_1_grant( bp_io_y_outChannels_2_credit_1_grant ),
       .io_outChannels_2_credit_0_grant( bp_io_y_outChannels_2_credit_0_grant ),
       .io_outChannels_1_flit_x( x_io_outChannels_1_flit_x ),
       .io_outChannels_1_flitValid( x_io_outChannels_1_flitValid ),
       .io_outChannels_1_credit_1_grant( bp_io_y_outChannels_1_credit_1_grant ),
       .io_outChannels_1_credit_0_grant( bp_io_y_outChannels_1_credit_0_grant ),
       .io_outChannels_0_flit_x( x_io_outChannels_0_flit_x ),
       .io_outChannels_0_flitValid( x_io_outChannels_0_flitValid ),
       .io_outChannels_0_credit_1_grant( bp_io_y_outChannels_0_credit_1_grant ),
       .io_outChannels_0_credit_0_grant( bp_io_y_outChannels_0_credit_0_grant ),
       //.io_counters_1_counterVal(  )
       //.io_counters_1_counterIndex(  )
       .io_counters_0_counterVal( x_io_counters_0_counterVal )
       //.io_counters_0_counterIndex(  )
       //.io_bypass(  )
  );
endmodule

module BusProbe_1(input clk, input reset,
    //input [54:0] io_inFlit_4_x
    //input [54:0] io_inFlit_3_x
    input [54:0] io_inFlit_2_x,
    input [54:0] io_inFlit_1_x,
    //input [54:0] io_inFlit_0_x
    input  io_inValid_4,
    input  io_inValid_3,
    input  io_inValid_2,
    input  io_inValid_1,
    input  io_inValid_0,
    input  io_routerCord,
    //input  io_startRecording
    output[15:0] io_cyclesChannelBusy_4,
    output[15:0] io_cyclesChannelBusy_3,
    output[15:0] io_cyclesChannelBusy_2,
    output[15:0] io_cyclesChannelBusy_1,
    output[15:0] io_cyclesChannelBusy_0,
    output[15:0] io_cyclesRouterBusy
);

  reg[0:0] T0;
  reg [15:0] cyclesRouterBusy;
  wire[15:0] T29;
  wire[15:0] T1;
  wire[15:0] T2;
  wire T3;
  wire[4:0] T4;
  wire[4:0] T5;
  wire[2:0] T6;
  wire[1:0] T7;
  reg  cyclesChannelBusyScoreboard_0;
  wire T30;
  wire T8;
  wire T9;
  reg  cyclesChannelBusyScoreboard_1;
  wire T31;
  wire T10;
  wire T11;
  reg  cyclesChannelBusyScoreboard_2;
  wire T32;
  wire T12;
  wire T13;
  wire[1:0] T14;
  reg  cyclesChannelBusyScoreboard_3;
  wire T33;
  wire T15;
  wire T16;
  reg  cyclesChannelBusyScoreboard_4;
  wire T34;
  wire T17;
  wire T18;
  reg [15:0] cyclesChannelBusy_0;
  wire[15:0] T35;
  wire[15:0] T19;
  wire[15:0] T20;
  reg [15:0] cyclesChannelBusy_1;
  wire[15:0] T36;
  wire[15:0] T21;
  wire[15:0] T22;
  reg [15:0] cyclesChannelBusy_2;
  wire[15:0] T37;
  wire[15:0] T23;
  wire[15:0] T24;
  reg [15:0] cyclesChannelBusy_3;
  wire[15:0] T38;
  wire[15:0] T25;
  wire[15:0] T26;
  reg [15:0] cyclesChannelBusy_4;
  wire[15:0] T39;
  wire[15:0] T27;
  wire[15:0] T28;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    T0 = 1'b0;
    cyclesRouterBusy = {1{1'b0}};
    cyclesChannelBusyScoreboard_0 = {1{1'b0}};
    cyclesChannelBusyScoreboard_1 = {1{1'b0}};
    cyclesChannelBusyScoreboard_2 = {1{1'b0}};
    cyclesChannelBusyScoreboard_3 = {1{1'b0}};
    cyclesChannelBusyScoreboard_4 = {1{1'b0}};
    cyclesChannelBusy_0 = {1{1'b0}};
    cyclesChannelBusy_1 = {1{1'b0}};
    cyclesChannelBusy_2 = {1{1'b0}};
    cyclesChannelBusy_3 = {1{1'b0}};
    cyclesChannelBusy_4 = {1{1'b0}};
  end
// synthesis translate_on
`endif

  assign io_cyclesRouterBusy = cyclesRouterBusy;
  assign T29 = reset ? 16'h0 : T1;
  assign T1 = T3 ? T2 : cyclesRouterBusy;
  assign T2 = cyclesRouterBusy + 16'h1;
  assign T3 = T4 != 5'h0;
  assign T4 = T5;
  assign T5 = {T14, T6};
  assign T6 = {cyclesChannelBusyScoreboard_2, T7};
  assign T7 = {cyclesChannelBusyScoreboard_1, cyclesChannelBusyScoreboard_0};
  assign T30 = reset ? 1'h0 : T8;
  assign T8 = T9 == 1'h0;
  assign T9 = io_inValid_0 ^ 1'h1;
  assign T31 = reset ? 1'h0 : T10;
  assign T10 = T11 == 1'h0;
  assign T11 = io_inValid_1 ^ 1'h1;
  assign T32 = reset ? 1'h0 : T12;
  assign T12 = T13 == 1'h0;
  assign T13 = io_inValid_2 ^ 1'h1;
  assign T14 = {cyclesChannelBusyScoreboard_4, cyclesChannelBusyScoreboard_3};
  assign T33 = reset ? 1'h0 : T15;
  assign T15 = T16 == 1'h0;
  assign T16 = io_inValid_3 ^ 1'h1;
  assign T34 = reset ? 1'h0 : T17;
  assign T17 = T18 == 1'h0;
  assign T18 = io_inValid_4 ^ 1'h1;
  assign io_cyclesChannelBusy_0 = cyclesChannelBusy_0;
  assign T35 = reset ? 16'h0 : T19;
  assign T19 = io_inValid_0 ? T20 : cyclesChannelBusy_0;
  assign T20 = cyclesChannelBusy_0 + 16'h1;
  assign io_cyclesChannelBusy_1 = cyclesChannelBusy_1;
  assign T36 = reset ? 16'h0 : T21;
  assign T21 = io_inValid_1 ? T22 : cyclesChannelBusy_1;
  assign T22 = cyclesChannelBusy_1 + 16'h1;
  assign io_cyclesChannelBusy_2 = cyclesChannelBusy_2;
  assign T37 = reset ? 16'h0 : T23;
  assign T23 = io_inValid_2 ? T24 : cyclesChannelBusy_2;
  assign T24 = cyclesChannelBusy_2 + 16'h1;
  assign io_cyclesChannelBusy_3 = cyclesChannelBusy_3;
  assign T38 = reset ? 16'h0 : T25;
  assign T25 = io_inValid_3 ? T26 : cyclesChannelBusy_3;
  assign T26 = cyclesChannelBusy_3 + 16'h1;
  assign io_cyclesChannelBusy_4 = cyclesChannelBusy_4;
  assign T39 = reset ? 16'h0 : T27;
  assign T27 = io_inValid_4 ? T28 : cyclesChannelBusy_4;
  assign T28 = cyclesChannelBusy_4 + 16'h1;

  always @(posedge clk) begin
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T0 <= 1'b1;
  if(!1'h1 && T0 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "BusProbe: RouterRadix must be > 1");
    $finish;
  end
// synthesis translate_on
`endif
    if(reset) begin
      cyclesRouterBusy <= 16'h0;
    end else if(T3) begin
      cyclesRouterBusy <= T2;
    end
    if(reset) begin
      cyclesChannelBusyScoreboard_0 <= 1'h0;
    end else begin
      cyclesChannelBusyScoreboard_0 <= T8;
    end
    if(reset) begin
      cyclesChannelBusyScoreboard_1 <= 1'h0;
    end else begin
      cyclesChannelBusyScoreboard_1 <= T10;
    end
    if(reset) begin
      cyclesChannelBusyScoreboard_2 <= 1'h0;
    end else begin
      cyclesChannelBusyScoreboard_2 <= T12;
    end
    if(reset) begin
      cyclesChannelBusyScoreboard_3 <= 1'h0;
    end else begin
      cyclesChannelBusyScoreboard_3 <= T15;
    end
    if(reset) begin
      cyclesChannelBusyScoreboard_4 <= 1'h0;
    end else begin
      cyclesChannelBusyScoreboard_4 <= T17;
    end
    if(reset) begin
      cyclesChannelBusy_0 <= 16'h0;
    end else if(io_inValid_0) begin
      cyclesChannelBusy_0 <= T20;
    end
    if(reset) begin
      cyclesChannelBusy_1 <= 16'h0;
    end else if(io_inValid_1) begin
      cyclesChannelBusy_1 <= T22;
    end
    if(reset) begin
      cyclesChannelBusy_2 <= 16'h0;
    end else if(io_inValid_2) begin
      cyclesChannelBusy_2 <= T24;
    end
    if(reset) begin
      cyclesChannelBusy_3 <= 16'h0;
    end else if(io_inValid_3) begin
      cyclesChannelBusy_3 <= T26;
    end
    if(reset) begin
      cyclesChannelBusy_4 <= 16'h0;
    end else if(io_inValid_4) begin
      cyclesChannelBusy_4 <= T28;
    end
  end
endmodule

module CMeshDOR_2(
    input [15:0] io_inHeadFlit_packetID,
    input  io_inHeadFlit_isTail,
    input  io_inHeadFlit_vcPort,
    input [3:0] io_inHeadFlit_packetType,
    input [1:0] io_inHeadFlit_destination_2,
    input [1:0] io_inHeadFlit_destination_1,
    input [1:0] io_inHeadFlit_destination_0,
    input [2:0] io_inHeadFlit_priorityLevel,
    output[15:0] io_outHeadFlit_packetID,
    output io_outHeadFlit_isTail,
    output io_outHeadFlit_vcPort,
    output[3:0] io_outHeadFlit_packetType,
    output[1:0] io_outHeadFlit_destination_2,
    output[1:0] io_outHeadFlit_destination_1,
    output[1:0] io_outHeadFlit_destination_0,
    output[2:0] io_outHeadFlit_priorityLevel,
    output[2:0] io_result,
    output[1:0] io_vcsAvailable_4,
    output[1:0] io_vcsAvailable_3,
    output[1:0] io_vcsAvailable_2,
    output[1:0] io_vcsAvailable_1,
    output[1:0] io_vcsAvailable_0
);

  wire[1:0] T0;
  wire[1:0] T26;
  wire T1;
  wire[1:0] T2;
  wire[1:0] T27;
  wire T3;
  wire[1:0] T4;
  wire[1:0] T28;
  wire T5;
  wire[1:0] T6;
  wire[1:0] T29;
  wire T7;
  wire[1:0] T8;
  wire[1:0] T30;
  wire T9;
  wire[2:0] T10;
  wire[2:0] resultReduction;
  wire[2:0] T11;
  wire[2:0] dimResults_1;
  wire[2:0] T12;
  wire[2:0] T31;
  wire[1:0] T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire[2:0] dimResults_0;
  wire[2:0] T32;
  wire[1:0] T18;
  wire[1:0] T33;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire[2:0] T34;
  wire T25;


  assign io_vcsAvailable_0 = T0;
  assign T0 = 2'h0 - T26;
  assign T26 = {1'h0, T1};
  assign T1 = io_result == 3'h0;
  assign io_vcsAvailable_1 = T2;
  assign T2 = 2'h0 - T27;
  assign T27 = {1'h0, T3};
  assign T3 = io_result == 3'h1;
  assign io_vcsAvailable_2 = T4;
  assign T4 = 2'h0 - T28;
  assign T28 = {1'h0, T5};
  assign T5 = io_result == 3'h2;
  assign io_vcsAvailable_3 = T6;
  assign T6 = 2'h0 - T29;
  assign T29 = {1'h0, T7};
  assign T7 = io_result == 3'h3;
  assign io_vcsAvailable_4 = T8;
  assign T8 = 2'h0 - T30;
  assign T30 = {1'h0, T9};
  assign T9 = io_result == 3'h4;
  assign io_result = T10;
  assign T10 = T25 ? T34 : resultReduction;
  assign resultReduction = T11;
  assign T11 = T24 ? dimResults_0 : dimResults_1;
  assign dimResults_1 = T12;
  assign T12 = T15 ? 3'h4 : T31;
  assign T31 = {1'h0, T13};
  assign T13 = T14 ? 2'h3 : 2'h0;
  assign T14 = 2'h0 < io_inHeadFlit_destination_1;
  assign T15 = T17 & T16;
  assign T16 = io_inHeadFlit_destination_1 < 2'h0;
  assign T17 = T14 ^ 1'h1;
  assign dimResults_0 = T32;
  assign T32 = {1'h0, T18};
  assign T18 = T21 ? 2'h2 : T33;
  assign T33 = {1'h0, T19};
  assign T19 = T20 ? 1'h1 : 1'h0;
  assign T20 = 2'h2 < io_inHeadFlit_destination_0;
  assign T21 = T23 & T22;
  assign T22 = io_inHeadFlit_destination_0 < 2'h2;
  assign T23 = T20 ^ 1'h1;
  assign T24 = dimResults_0 != 3'h0;
  assign T34 = {1'h0, io_inHeadFlit_destination_2};
  assign T25 = resultReduction == 3'h0;
  assign io_outHeadFlit_priorityLevel = io_inHeadFlit_priorityLevel;
  assign io_outHeadFlit_destination_0 = io_inHeadFlit_destination_0;
  assign io_outHeadFlit_destination_1 = io_inHeadFlit_destination_1;
  assign io_outHeadFlit_destination_2 = io_inHeadFlit_destination_2;
  assign io_outHeadFlit_packetType = io_inHeadFlit_packetType;
  assign io_outHeadFlit_vcPort = io_inHeadFlit_vcPort;
  assign io_outHeadFlit_isTail = io_inHeadFlit_isTail;
  assign io_outHeadFlit_packetID = io_inHeadFlit_packetID;
endmodule

module SimpleVCRouter_2((* gated_clock = "true" *) input clk, input reset,
    input [54:0] io_inChannels_4_flit_x,
    input  io_inChannels_4_flitValid,
    output io_inChannels_4_credit_1_grant,
    output io_inChannels_4_credit_0_grant,
    input [54:0] io_inChannels_3_flit_x,
    input  io_inChannels_3_flitValid,
    output io_inChannels_3_credit_1_grant,
    output io_inChannels_3_credit_0_grant,
    input [54:0] io_inChannels_2_flit_x,
    input  io_inChannels_2_flitValid,
    output io_inChannels_2_credit_1_grant,
    output io_inChannels_2_credit_0_grant,
    input [54:0] io_inChannels_1_flit_x,
    input  io_inChannels_1_flitValid,
    output io_inChannels_1_credit_1_grant,
    output io_inChannels_1_credit_0_grant,
    input [54:0] io_inChannels_0_flit_x,
    input  io_inChannels_0_flitValid,
    output io_inChannels_0_credit_1_grant,
    output io_inChannels_0_credit_0_grant,
    output[54:0] io_outChannels_4_flit_x,
    output io_outChannels_4_flitValid,
    input  io_outChannels_4_credit_1_grant,
    input  io_outChannels_4_credit_0_grant,
    output[54:0] io_outChannels_3_flit_x,
    output io_outChannels_3_flitValid,
    input  io_outChannels_3_credit_1_grant,
    input  io_outChannels_3_credit_0_grant,
    output[54:0] io_outChannels_2_flit_x,
    output io_outChannels_2_flitValid,
    input  io_outChannels_2_credit_1_grant,
    input  io_outChannels_2_credit_0_grant,
    output[54:0] io_outChannels_1_flit_x,
    output io_outChannels_1_flitValid,
    input  io_outChannels_1_credit_1_grant,
    input  io_outChannels_1_credit_0_grant,
    output[54:0] io_outChannels_0_flit_x,
    output io_outChannels_0_flitValid,
    input  io_outChannels_0_credit_1_grant,
    input  io_outChannels_0_credit_0_grant,
    //output[31:0] io_counters_1_counterVal
    //output[7:0] io_counters_1_counterIndex
    output[31:0] io_counters_0_counterVal
    //output[7:0] io_counters_0_counterIndex
    //input  io_bypass
);

  reg[0:0] T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  wire[53:0] T8;
  wire T9;
  wire[30:0] T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  reg[0:0] T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  reg[0:0] T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire[53:0] T30;
  wire T31;
  wire[30:0] T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  reg[0:0] T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  reg[0:0] T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire[53:0] T52;
  wire T53;
  wire[30:0] T54;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  reg[0:0] T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  reg[0:0] T66;
  wire T67;
  wire T68;
  wire T69;
  wire T70;
  wire T71;
  wire T72;
  wire T73;
  wire[53:0] T74;
  wire T75;
  wire[30:0] T76;
  wire T77;
  wire T78;
  wire T79;
  wire T80;
  wire T81;
  wire T82;
  reg[0:0] T83;
  wire T84;
  wire T85;
  wire T86;
  wire T87;
  reg[0:0] T88;
  wire T89;
  wire T90;
  wire T91;
  wire T92;
  wire T93;
  wire T94;
  wire T95;
  wire[53:0] T96;
  wire T97;
  wire[30:0] T98;
  wire T99;
  wire T100;
  wire T101;
  wire T102;
  wire T103;
  wire T104;
  reg[0:0] T105;
  wire T106;
  wire T107;
  wire T108;
  wire T109;
  reg[0:0] T110;
  wire T111;
  wire T112;
  wire T113;
  wire T114;
  wire T115;
  wire T116;
  wire T117;
  wire[53:0] T118;
  wire T119;
  wire[30:0] T120;
  wire T121;
  wire T122;
  wire T123;
  wire T124;
  wire T125;
  wire T126;
  reg[0:0] T127;
  wire T128;
  wire T129;
  wire T130;
  wire T131;
  reg[0:0] T132;
  wire T133;
  wire T134;
  wire T135;
  wire T136;
  wire T137;
  wire T138;
  wire T139;
  wire[53:0] T140;
  wire T141;
  wire[30:0] T142;
  wire T143;
  wire T144;
  wire T145;
  wire T146;
  wire T147;
  wire T148;
  reg[0:0] T149;
  wire T150;
  wire T151;
  wire T152;
  wire T153;
  reg[0:0] T154;
  wire T155;
  wire T156;
  wire T157;
  wire T158;
  wire T159;
  wire T160;
  wire T161;
  wire[53:0] T162;
  wire T163;
  wire[30:0] T164;
  wire T165;
  wire T166;
  wire T167;
  wire T168;
  wire T169;
  wire T170;
  reg[0:0] T171;
  wire T172;
  wire T173;
  wire T174;
  wire T175;
  reg[0:0] T176;
  wire T177;
  wire T178;
  wire T179;
  wire T180;
  wire T181;
  wire T182;
  wire T183;
  wire[53:0] T184;
  wire T185;
  wire[30:0] T186;
  wire T187;
  wire T188;
  wire T189;
  wire T190;
  wire T191;
  wire T192;
  reg[0:0] T193;
  wire T194;
  wire T195;
  wire T196;
  wire T197;
  reg[0:0] T198;
  wire T199;
  wire T200;
  wire T201;
  wire T202;
  wire T203;
  wire T204;
  wire T205;
  wire[53:0] T206;
  wire T207;
  wire[30:0] T208;
  wire T209;
  wire T210;
  wire T211;
  wire T212;
  wire T213;
  wire T214;
  reg[0:0] T215;
  wire T216;
  wire T217;
  wire T218;
  wire T219;
  wire T220;
  wire T221;
  wire T222;
  wire T223;
  wire T224;
  wire[53:0] T225;
  wire T226;
  wire[30:0] T227;
  wire T228;
  wire T229;
  wire T230;
  wire T231;
  wire T232;
  wire T233;
  wire T234;
  wire T235;
  wire T236;
  wire[53:0] T237;
  wire T238;
  wire[30:0] T239;
  wire T240;
  wire T241;
  wire T242;
  wire T243;
  wire T244;
  wire T245;
  wire T246;
  wire T247;
  wire T248;
  wire[53:0] T249;
  wire T250;
  wire[30:0] T251;
  wire T252;
  wire T253;
  wire T254;
  wire T255;
  wire T256;
  wire T257;
  wire T258;
  wire T259;
  wire T260;
  wire[53:0] T261;
  wire T262;
  wire[30:0] T263;
  wire T264;
  wire T265;
  wire T266;
  wire T267;
  wire T268;
  wire T269;
  wire T270;
  wire T271;
  wire T272;
  wire[53:0] T273;
  wire T274;
  wire[30:0] T275;
  wire T276;
  wire T277;
  wire T278;
  wire T279;
  wire[54:0] T280;
  wire[54:0] T281;
  wire T3112;
  reg [54:0] R282;
  wire[54:0] T3113;
  wire[54:0] T283;
  wire[54:0] T3114;
  wire T284;
  wire T285;
  wire[54:0] T286;
  wire[54:0] T287;
  wire T288;
  wire T289;
  wire[1:0] T290;
  wire[1:0] T291;
  wire[1:0] T292;
  wire T293;
  wire[2:0] T294;
  reg [2:0] R295;
  wire[2:0] T3115;
  wire[1:0] T296;
  wire T297;
  wire T298;
  wire T299;
  wire T300;
  wire T301;
  wire T302;
  wire T303;
  wire T304;
  wire creditConsReady_0_0;
  wire creditConsReady_1_0;
  wire T305;
  wire[2:0] T306;
  wire T307;
  wire creditConsReady_2_0;
  wire creditConsReady_3_0;
  wire T308;
  wire T309;
  wire creditConsReady_4_0;
  wire T310;
  wire T311;
  wire T312;
  wire T313;
  wire creditConsReady_0_1;
  wire creditConsReady_1_1;
  wire T314;
  wire T315;
  wire creditConsReady_2_1;
  wire creditConsReady_3_1;
  wire T316;
  wire T317;
  wire creditConsReady_4_1;
  wire T318;
  wire T319;
  wire T3116;
  wire T320;
  wire T321;
  wire[3:0] T322;
  wire[3:0] T323;
  wire[3:0] T324;
  wire T325;
  wire[2:0] T326;
  wire[3:0] T327;
  wire T328;
  wire T329;
  wire T330;
  wire T331;
  wire T332;
  wire T333;
  wire T334;
  wire[2:0] T335;
  wire T336;
  wire T337;
  wire T338;
  wire T339;
  wire T340;
  wire T341;
  wire T342;
  wire T343;
  wire[53:0] T344;
  wire T345;
  wire[30:0] T346;
  wire T347;
  wire T348;
  reg  R349;
  wire T3117;
  wire[2:0] T350;
  wire[30:0] T351;
  wire[54:0] T352;
  wire[1:0] T353;
  wire[1:0] T354;
  wire[1:0] T355;
  wire[3:0] T356;
  wire T357;
  wire T358;
  wire[15:0] T359;
  wire T360;
  wire T361;
  wire T362;
  wire T363;
  wire T364;
  wire T365;
  wire T366;
  wire T367;
  wire T368;
  wire T369;
  wire T370;
  wire T371;
  wire T372;
  wire T373;
  wire T374;
  wire T375;
  wire T376;
  wire T377;
  wire T378;
  wire T379;
  wire T380;
  wire T381;
  wire T382;
  wire T383;
  wire T384;
  wire T385;
  wire T386;
  wire T387;
  wire[54:0] T3118;
  wire[30:0] T388;
  wire[30:0] T389;
  wire[8:0] T390;
  wire[4:0] T391;
  wire[3:0] T392;
  wire[21:0] T393;
  wire[4:0] T394;
  wire[16:0] T395;
  wire T396;
  wire T397;
  wire T398;
  wire T399;
  wire flitsAreTail_9;
  wire T400;
  wire T401;
  wire T402;
  wire T403;
  wire[53:0] T404;
  wire T405;
  wire[30:0] T406;
  wire T407;
  wire T408;
  wire T409;
  wire T410;
  wire T411;
  wire[54:0] T412;
  wire[54:0] T413;
  wire T414;
  wire T415;
  wire T416;
  wire T417;
  wire T418;
  wire T419;
  wire T420;
  wire T421;
  wire T422;
  wire T423;
  wire[54:0] T424;
  wire[54:0] T425;
  wire T3119;
  reg [54:0] R426;
  wire[54:0] T3120;
  wire[54:0] T427;
  wire[54:0] T3121;
  wire T428;
  wire T429;
  wire[54:0] T430;
  wire[54:0] T431;
  wire T432;
  wire T433;
  wire[1:0] T434;
  wire[1:0] T435;
  wire[1:0] T436;
  wire T437;
  wire[2:0] T438;
  reg [2:0] R439;
  wire[2:0] T3122;
  wire[1:0] T440;
  wire T441;
  wire T442;
  wire T443;
  wire T444;
  wire T445;
  wire T446;
  wire T447;
  wire T448;
  wire T449;
  wire[2:0] T450;
  wire T451;
  wire T452;
  wire T453;
  wire T454;
  wire T455;
  wire T456;
  wire T457;
  wire T458;
  wire T459;
  wire T460;
  wire T461;
  wire T462;
  wire T463;
  wire T3123;
  wire T464;
  wire T465;
  wire[3:0] T466;
  wire[3:0] T467;
  wire[3:0] T468;
  wire T469;
  wire[2:0] T470;
  wire[3:0] T471;
  wire T472;
  wire T473;
  wire T474;
  wire T475;
  wire T476;
  wire T477;
  wire T478;
  wire[2:0] T479;
  wire T480;
  wire T481;
  wire T482;
  wire T483;
  wire T484;
  wire T485;
  wire T486;
  wire T487;
  wire[53:0] T488;
  wire T489;
  wire[30:0] T490;
  wire T491;
  wire T492;
  reg  R493;
  wire T3124;
  wire[2:0] T494;
  wire[30:0] T495;
  wire[54:0] T496;
  wire[1:0] T497;
  wire[1:0] T498;
  wire[1:0] T499;
  wire[3:0] T500;
  wire T501;
  wire T502;
  wire[15:0] T503;
  wire T504;
  wire T505;
  wire T506;
  wire T507;
  wire T508;
  wire T509;
  wire T510;
  wire T511;
  wire T512;
  wire T513;
  wire T514;
  wire T515;
  wire T516;
  wire T517;
  wire T518;
  wire T519;
  wire T520;
  wire T521;
  wire T522;
  wire T523;
  wire T524;
  wire T525;
  wire T526;
  wire T527;
  wire T528;
  wire T529;
  wire T530;
  wire T531;
  wire[54:0] T3125;
  wire[30:0] T532;
  wire[30:0] T533;
  wire[8:0] T534;
  wire[4:0] T535;
  wire[3:0] T536;
  wire[21:0] T537;
  wire[4:0] T538;
  wire[16:0] T539;
  wire T540;
  wire T541;
  wire T542;
  wire T543;
  wire flitsAreTail_8;
  wire T544;
  wire T545;
  wire T546;
  wire T547;
  wire[53:0] T548;
  wire T549;
  wire[30:0] T550;
  wire T551;
  wire T552;
  wire T553;
  wire T554;
  wire T555;
  wire[54:0] T556;
  wire[54:0] T557;
  wire T558;
  wire T559;
  wire T560;
  wire T561;
  wire T562;
  wire T563;
  wire T564;
  wire T565;
  wire T566;
  wire T567;
  wire[54:0] T568;
  wire[54:0] T569;
  wire T3126;
  reg [54:0] R570;
  wire[54:0] T3127;
  wire[54:0] T571;
  wire[54:0] T3128;
  wire T572;
  wire T573;
  wire[54:0] T574;
  wire[54:0] T575;
  wire T576;
  wire T577;
  wire[1:0] T578;
  wire[1:0] T579;
  wire[1:0] T580;
  wire T581;
  wire[2:0] T582;
  reg [2:0] R583;
  wire[2:0] T3129;
  wire[1:0] T584;
  wire T585;
  wire T586;
  wire T587;
  wire T588;
  wire T589;
  wire T590;
  wire T591;
  wire T592;
  wire T593;
  wire[2:0] T594;
  wire T595;
  wire T596;
  wire T597;
  wire T598;
  wire T599;
  wire T600;
  wire T601;
  wire T602;
  wire T603;
  wire T604;
  wire T605;
  wire T606;
  wire T607;
  wire T3130;
  wire T608;
  wire T609;
  wire[3:0] T610;
  wire[3:0] T611;
  wire[3:0] T612;
  wire T613;
  wire[2:0] T614;
  wire[3:0] T615;
  wire T616;
  wire T617;
  wire T618;
  wire T619;
  wire T620;
  wire T621;
  wire T622;
  wire[2:0] T623;
  wire T624;
  wire T625;
  wire T626;
  wire T627;
  wire T628;
  wire T629;
  wire T630;
  wire T631;
  wire[53:0] T632;
  wire T633;
  wire[30:0] T634;
  wire T635;
  wire T636;
  reg  R637;
  wire T3131;
  wire[2:0] T638;
  wire[30:0] T639;
  wire[54:0] T640;
  wire[1:0] T641;
  wire[1:0] T642;
  wire[1:0] T643;
  wire[3:0] T644;
  wire T645;
  wire T646;
  wire[15:0] T647;
  wire T648;
  wire T649;
  wire T650;
  wire T651;
  wire T652;
  wire T653;
  wire T654;
  wire T655;
  wire T656;
  wire T657;
  wire T658;
  wire T659;
  wire T660;
  wire T661;
  wire T662;
  wire T663;
  wire T664;
  wire T665;
  wire T666;
  wire T667;
  wire T668;
  wire T669;
  wire T670;
  wire T671;
  wire T672;
  wire T673;
  wire T674;
  wire T675;
  wire[54:0] T3132;
  wire[30:0] T676;
  wire[30:0] T677;
  wire[8:0] T678;
  wire[4:0] T679;
  wire[3:0] T680;
  wire[21:0] T681;
  wire[4:0] T682;
  wire[16:0] T683;
  wire T684;
  wire T685;
  wire T686;
  wire T687;
  wire flitsAreTail_7;
  wire T688;
  wire T689;
  wire T690;
  wire T691;
  wire[53:0] T692;
  wire T693;
  wire[30:0] T694;
  wire T695;
  wire T696;
  wire T697;
  wire T698;
  wire T699;
  wire[54:0] T700;
  wire[54:0] T701;
  wire T702;
  wire T703;
  wire T704;
  wire T705;
  wire T706;
  wire T707;
  wire T708;
  wire T709;
  wire T710;
  wire T711;
  wire[54:0] T712;
  wire[54:0] T713;
  wire T3133;
  reg [54:0] R714;
  wire[54:0] T3134;
  wire[54:0] T715;
  wire[54:0] T3135;
  wire T716;
  wire T717;
  wire[54:0] T718;
  wire[54:0] T719;
  wire T720;
  wire T721;
  wire[1:0] T722;
  wire[1:0] T723;
  wire[1:0] T724;
  wire T725;
  wire[2:0] T726;
  reg [2:0] R727;
  wire[2:0] T3136;
  wire[1:0] T728;
  wire T729;
  wire T730;
  wire T731;
  wire T732;
  wire T733;
  wire T734;
  wire T735;
  wire T736;
  wire T737;
  wire[2:0] T738;
  wire T739;
  wire T740;
  wire T741;
  wire T742;
  wire T743;
  wire T744;
  wire T745;
  wire T746;
  wire T747;
  wire T748;
  wire T749;
  wire T750;
  wire T751;
  wire T3137;
  wire T752;
  wire T753;
  wire[3:0] T754;
  wire[3:0] T755;
  wire[3:0] T756;
  wire T757;
  wire[2:0] T758;
  wire[3:0] T759;
  wire T760;
  wire T761;
  wire T762;
  wire T763;
  wire T764;
  wire T765;
  wire T766;
  wire[2:0] T767;
  wire T768;
  wire T769;
  wire T770;
  wire T771;
  wire T772;
  wire T773;
  wire T774;
  wire T775;
  wire[53:0] T776;
  wire T777;
  wire[30:0] T778;
  wire T779;
  wire T780;
  reg  R781;
  wire T3138;
  wire[2:0] T782;
  wire[30:0] T783;
  wire[54:0] T784;
  wire[1:0] T785;
  wire[1:0] T786;
  wire[1:0] T787;
  wire[3:0] T788;
  wire T789;
  wire T790;
  wire[15:0] T791;
  wire T792;
  wire T793;
  wire T794;
  wire T795;
  wire T796;
  wire T797;
  wire T798;
  wire T799;
  wire T800;
  wire T801;
  wire T802;
  wire T803;
  wire T804;
  wire T805;
  wire T806;
  wire T807;
  wire T808;
  wire T809;
  wire T810;
  wire T811;
  wire T812;
  wire T813;
  wire T814;
  wire T815;
  wire T816;
  wire T817;
  wire T818;
  wire T819;
  wire[54:0] T3139;
  wire[30:0] T820;
  wire[30:0] T821;
  wire[8:0] T822;
  wire[4:0] T823;
  wire[3:0] T824;
  wire[21:0] T825;
  wire[4:0] T826;
  wire[16:0] T827;
  wire T828;
  wire T829;
  wire T830;
  wire T831;
  wire flitsAreTail_6;
  wire T832;
  wire T833;
  wire T834;
  wire T835;
  wire[53:0] T836;
  wire T837;
  wire[30:0] T838;
  wire T839;
  wire T840;
  wire T841;
  wire T842;
  wire T843;
  wire[54:0] T844;
  wire[54:0] T845;
  wire T846;
  wire T847;
  wire T848;
  wire T849;
  wire T850;
  wire T851;
  wire T852;
  wire T853;
  wire T854;
  wire T855;
  wire[54:0] T856;
  wire[54:0] T857;
  wire T3140;
  reg [54:0] R858;
  wire[54:0] T3141;
  wire[54:0] T859;
  wire[54:0] T3142;
  wire T860;
  wire T861;
  wire[54:0] T862;
  wire[54:0] T863;
  wire T864;
  wire T865;
  wire[1:0] T866;
  wire[1:0] T867;
  wire[1:0] T868;
  wire T869;
  wire[2:0] T870;
  reg [2:0] R871;
  wire[2:0] T3143;
  wire[1:0] T872;
  wire T873;
  wire T874;
  wire T875;
  wire T876;
  wire T877;
  wire T878;
  wire T879;
  wire T880;
  wire T881;
  wire[2:0] T882;
  wire T883;
  wire T884;
  wire T885;
  wire T886;
  wire T887;
  wire T888;
  wire T889;
  wire T890;
  wire T891;
  wire T892;
  wire T893;
  wire T894;
  wire T895;
  wire T3144;
  wire T896;
  wire T897;
  wire[3:0] T898;
  wire[3:0] T899;
  wire[3:0] T900;
  wire T901;
  wire[2:0] T902;
  wire[3:0] T903;
  wire T904;
  wire T905;
  wire T906;
  wire T907;
  wire T908;
  wire T909;
  wire T910;
  wire[2:0] T911;
  wire T912;
  wire T913;
  wire T914;
  wire T915;
  wire T916;
  wire T917;
  wire T918;
  wire T919;
  wire[53:0] T920;
  wire T921;
  wire[30:0] T922;
  wire T923;
  wire T924;
  reg  R925;
  wire T3145;
  wire[2:0] T926;
  wire[30:0] T927;
  wire[54:0] T928;
  wire[1:0] T929;
  wire[1:0] T930;
  wire[1:0] T931;
  wire[3:0] T932;
  wire T933;
  wire T934;
  wire[15:0] T935;
  wire T936;
  wire T937;
  wire T938;
  wire T939;
  wire T940;
  wire T941;
  wire T942;
  wire T943;
  wire T944;
  wire T945;
  wire T946;
  wire T947;
  wire T948;
  wire T949;
  wire T950;
  wire T951;
  wire T952;
  wire T953;
  wire T954;
  wire T955;
  wire T956;
  wire T957;
  wire T958;
  wire T959;
  wire T960;
  wire T961;
  wire T962;
  wire T963;
  wire[54:0] T3146;
  wire[30:0] T964;
  wire[30:0] T965;
  wire[8:0] T966;
  wire[4:0] T967;
  wire[3:0] T968;
  wire[21:0] T969;
  wire[4:0] T970;
  wire[16:0] T971;
  wire T972;
  wire T973;
  wire T974;
  wire T975;
  wire flitsAreTail_5;
  wire T976;
  wire T977;
  wire T978;
  wire T979;
  wire[53:0] T980;
  wire T981;
  wire[30:0] T982;
  wire T983;
  wire T984;
  wire T985;
  wire T986;
  wire T987;
  wire[54:0] T988;
  wire[54:0] T989;
  wire T990;
  wire T991;
  wire T992;
  wire T993;
  wire T994;
  wire T995;
  wire T996;
  wire T997;
  wire T998;
  wire T999;
  wire[54:0] T1000;
  wire[54:0] T1001;
  wire T3147;
  reg [54:0] R1002;
  wire[54:0] T3148;
  wire[54:0] T1003;
  wire[54:0] T3149;
  wire T1004;
  wire T1005;
  wire[54:0] T1006;
  wire[54:0] T1007;
  wire T1008;
  wire T1009;
  wire[1:0] T1010;
  wire[1:0] T1011;
  wire[1:0] T1012;
  wire T1013;
  wire[2:0] T1014;
  reg [2:0] R1015;
  wire[2:0] T3150;
  wire[1:0] T1016;
  wire T1017;
  wire T1018;
  wire T1019;
  wire T1020;
  wire T1021;
  wire T1022;
  wire T1023;
  wire T1024;
  wire T1025;
  wire[2:0] T1026;
  wire T1027;
  wire T1028;
  wire T1029;
  wire T1030;
  wire T1031;
  wire T1032;
  wire T1033;
  wire T1034;
  wire T1035;
  wire T1036;
  wire T1037;
  wire T1038;
  wire T1039;
  wire T3151;
  wire T1040;
  wire T1041;
  wire[3:0] T1042;
  wire[3:0] T1043;
  wire[3:0] T1044;
  wire T1045;
  wire[2:0] T1046;
  wire[3:0] T1047;
  wire T1048;
  wire T1049;
  wire T1050;
  wire T1051;
  wire T1052;
  wire T1053;
  wire T1054;
  wire[2:0] T1055;
  wire T1056;
  wire T1057;
  wire T1058;
  wire T1059;
  wire T1060;
  wire T1061;
  wire T1062;
  wire T1063;
  wire[53:0] T1064;
  wire T1065;
  wire[30:0] T1066;
  wire T1067;
  wire T1068;
  reg  R1069;
  wire T3152;
  wire[2:0] T1070;
  wire[30:0] T1071;
  wire[54:0] T1072;
  wire[1:0] T1073;
  wire[1:0] T1074;
  wire[1:0] T1075;
  wire[3:0] T1076;
  wire T1077;
  wire T1078;
  wire[15:0] T1079;
  wire T1080;
  wire T1081;
  wire T1082;
  wire T1083;
  wire T1084;
  wire T1085;
  wire T1086;
  wire T1087;
  wire T1088;
  wire T1089;
  wire T1090;
  wire T1091;
  wire T1092;
  wire T1093;
  wire T1094;
  wire T1095;
  wire T1096;
  wire T1097;
  wire T1098;
  wire T1099;
  wire T1100;
  wire T1101;
  wire T1102;
  wire T1103;
  wire T1104;
  wire T1105;
  wire T1106;
  wire T1107;
  wire[54:0] T3153;
  wire[30:0] T1108;
  wire[30:0] T1109;
  wire[8:0] T1110;
  wire[4:0] T1111;
  wire[3:0] T1112;
  wire[21:0] T1113;
  wire[4:0] T1114;
  wire[16:0] T1115;
  wire T1116;
  wire T1117;
  wire T1118;
  wire T1119;
  wire flitsAreTail_4;
  wire T1120;
  wire T1121;
  wire T1122;
  wire T1123;
  wire[53:0] T1124;
  wire T1125;
  wire[30:0] T1126;
  wire T1127;
  wire T1128;
  wire T1129;
  wire T1130;
  wire T1131;
  wire[54:0] T1132;
  wire[54:0] T1133;
  wire T1134;
  wire T1135;
  wire T1136;
  wire T1137;
  wire T1138;
  wire T1139;
  wire T1140;
  wire T1141;
  wire T1142;
  wire T1143;
  wire[54:0] T1144;
  wire[54:0] T1145;
  wire T3154;
  reg [54:0] R1146;
  wire[54:0] T3155;
  wire[54:0] T1147;
  wire[54:0] T3156;
  wire T1148;
  wire T1149;
  wire[54:0] T1150;
  wire[54:0] T1151;
  wire T1152;
  wire T1153;
  wire[1:0] T1154;
  wire[1:0] T1155;
  wire[1:0] T1156;
  wire T1157;
  wire[2:0] T1158;
  reg [2:0] R1159;
  wire[2:0] T3157;
  wire[1:0] T1160;
  wire T1161;
  wire T1162;
  wire T1163;
  wire T1164;
  wire T1165;
  wire T1166;
  wire T1167;
  wire T1168;
  wire T1169;
  wire[2:0] T1170;
  wire T1171;
  wire T1172;
  wire T1173;
  wire T1174;
  wire T1175;
  wire T1176;
  wire T1177;
  wire T1178;
  wire T1179;
  wire T1180;
  wire T1181;
  wire T1182;
  wire T1183;
  wire T3158;
  wire T1184;
  wire T1185;
  wire[3:0] T1186;
  wire[3:0] T1187;
  wire[3:0] T1188;
  wire T1189;
  wire[2:0] T1190;
  wire[3:0] T1191;
  wire T1192;
  wire T1193;
  wire T1194;
  wire T1195;
  wire T1196;
  wire T1197;
  wire T1198;
  wire[2:0] T1199;
  wire T1200;
  wire T1201;
  wire T1202;
  wire T1203;
  wire T1204;
  wire T1205;
  wire T1206;
  wire T1207;
  wire[53:0] T1208;
  wire T1209;
  wire[30:0] T1210;
  wire T1211;
  wire T1212;
  reg  R1213;
  wire T3159;
  wire[2:0] T1214;
  wire[30:0] T1215;
  wire[54:0] T1216;
  wire[1:0] T1217;
  wire[1:0] T1218;
  wire[1:0] T1219;
  wire[3:0] T1220;
  wire T1221;
  wire T1222;
  wire[15:0] T1223;
  wire T1224;
  wire T1225;
  wire T1226;
  wire T1227;
  wire T1228;
  wire T1229;
  wire T1230;
  wire T1231;
  wire T1232;
  wire T1233;
  wire T1234;
  wire T1235;
  wire T1236;
  wire T1237;
  wire T1238;
  wire T1239;
  wire T1240;
  wire T1241;
  wire T1242;
  wire T1243;
  wire T1244;
  wire T1245;
  wire T1246;
  wire T1247;
  wire T1248;
  wire T1249;
  wire T1250;
  wire T1251;
  wire[54:0] T3160;
  wire[30:0] T1252;
  wire[30:0] T1253;
  wire[8:0] T1254;
  wire[4:0] T1255;
  wire[3:0] T1256;
  wire[21:0] T1257;
  wire[4:0] T1258;
  wire[16:0] T1259;
  wire T1260;
  wire T1261;
  wire T1262;
  wire T1263;
  wire flitsAreTail_3;
  wire T1264;
  wire T1265;
  wire T1266;
  wire T1267;
  wire[53:0] T1268;
  wire T1269;
  wire[30:0] T1270;
  wire T1271;
  wire T1272;
  wire T1273;
  wire T1274;
  wire T1275;
  wire[54:0] T1276;
  wire[54:0] T1277;
  wire T1278;
  wire T1279;
  wire T1280;
  wire T1281;
  wire T1282;
  wire T1283;
  wire T1284;
  wire T1285;
  wire T1286;
  wire T1287;
  wire[54:0] T1288;
  wire[54:0] T1289;
  wire T3161;
  reg [54:0] R1290;
  wire[54:0] T3162;
  wire[54:0] T1291;
  wire[54:0] T3163;
  wire T1292;
  wire T1293;
  wire[54:0] T1294;
  wire[54:0] T1295;
  wire T1296;
  wire T1297;
  wire[1:0] T1298;
  wire[1:0] T1299;
  wire[1:0] T1300;
  wire T1301;
  wire[2:0] T1302;
  reg [2:0] R1303;
  wire[2:0] T3164;
  wire[1:0] T1304;
  wire T1305;
  wire T1306;
  wire T1307;
  wire T1308;
  wire T1309;
  wire T1310;
  wire T1311;
  wire T1312;
  wire T1313;
  wire[2:0] T1314;
  wire T1315;
  wire T1316;
  wire T1317;
  wire T1318;
  wire T1319;
  wire T1320;
  wire T1321;
  wire T1322;
  wire T1323;
  wire T1324;
  wire T1325;
  wire T1326;
  wire T1327;
  wire T3165;
  wire T1328;
  wire T1329;
  wire[3:0] T1330;
  wire[3:0] T1331;
  wire[3:0] T1332;
  wire T1333;
  wire[2:0] T1334;
  wire[3:0] T1335;
  wire T1336;
  wire T1337;
  wire T1338;
  wire T1339;
  wire T1340;
  wire T1341;
  wire T1342;
  wire[2:0] T1343;
  wire T1344;
  wire T1345;
  wire T1346;
  wire T1347;
  wire T1348;
  wire T1349;
  wire T1350;
  wire T1351;
  wire[53:0] T1352;
  wire T1353;
  wire[30:0] T1354;
  wire T1355;
  wire T1356;
  reg  R1357;
  wire T3166;
  wire[2:0] T1358;
  wire[30:0] T1359;
  wire[54:0] T1360;
  wire[1:0] T1361;
  wire[1:0] T1362;
  wire[1:0] T1363;
  wire[3:0] T1364;
  wire T1365;
  wire T1366;
  wire[15:0] T1367;
  wire T1368;
  wire T1369;
  wire T1370;
  wire T1371;
  wire T1372;
  wire T1373;
  wire T1374;
  wire T1375;
  wire T1376;
  wire T1377;
  wire T1378;
  wire T1379;
  wire T1380;
  wire T1381;
  wire T1382;
  wire T1383;
  wire T1384;
  wire T1385;
  wire T1386;
  wire T1387;
  wire T1388;
  wire T1389;
  wire T1390;
  wire T1391;
  wire T1392;
  wire T1393;
  wire T1394;
  wire T1395;
  wire[54:0] T3167;
  wire[30:0] T1396;
  wire[30:0] T1397;
  wire[8:0] T1398;
  wire[4:0] T1399;
  wire[3:0] T1400;
  wire[21:0] T1401;
  wire[4:0] T1402;
  wire[16:0] T1403;
  wire T1404;
  wire T1405;
  wire T1406;
  wire T1407;
  wire flitsAreTail_2;
  wire T1408;
  wire T1409;
  wire T1410;
  wire T1411;
  wire[53:0] T1412;
  wire T1413;
  wire[30:0] T1414;
  wire T1415;
  wire T1416;
  wire T1417;
  wire T1418;
  wire T1419;
  wire[54:0] T1420;
  wire[54:0] T1421;
  wire T1422;
  wire T1423;
  wire T1424;
  wire T1425;
  wire T1426;
  wire T1427;
  wire T1428;
  wire T1429;
  wire T1430;
  wire T1431;
  wire[54:0] T1432;
  wire[54:0] T1433;
  wire T3168;
  reg [54:0] R1434;
  wire[54:0] T3169;
  wire[54:0] T1435;
  wire[54:0] T3170;
  wire T1436;
  wire T1437;
  wire[54:0] T1438;
  wire[54:0] T1439;
  wire T1440;
  wire T1441;
  wire[1:0] T1442;
  wire[1:0] T1443;
  wire[1:0] T1444;
  wire T1445;
  wire[2:0] T1446;
  reg [2:0] R1447;
  wire[2:0] T3171;
  wire[1:0] T1448;
  wire T1449;
  wire T1450;
  wire T1451;
  wire T1452;
  wire T1453;
  wire T1454;
  wire T1455;
  wire T1456;
  wire T1457;
  wire[2:0] T1458;
  wire T1459;
  wire T1460;
  wire T1461;
  wire T1462;
  wire T1463;
  wire T1464;
  wire T1465;
  wire T1466;
  wire T1467;
  wire T1468;
  wire T1469;
  wire T1470;
  wire T1471;
  wire T3172;
  wire T1472;
  wire T1473;
  wire[3:0] T1474;
  wire[3:0] T1475;
  wire[3:0] T1476;
  wire T1477;
  wire[2:0] T1478;
  wire[3:0] T1479;
  wire T1480;
  wire T1481;
  wire T1482;
  wire T1483;
  wire T1484;
  wire T1485;
  wire T1486;
  wire[2:0] T1487;
  wire T1488;
  wire T1489;
  wire T1490;
  wire T1491;
  wire T1492;
  wire T1493;
  wire T1494;
  wire T1495;
  wire[53:0] T1496;
  wire T1497;
  wire[30:0] T1498;
  wire T1499;
  wire T1500;
  reg  R1501;
  wire T3173;
  wire[2:0] T1502;
  wire[30:0] T1503;
  wire[54:0] T1504;
  wire[1:0] T1505;
  wire[1:0] T1506;
  wire[1:0] T1507;
  wire[3:0] T1508;
  wire T1509;
  wire T1510;
  wire[15:0] T1511;
  wire T1512;
  wire T1513;
  wire T1514;
  wire T1515;
  wire T1516;
  wire T1517;
  wire T1518;
  wire T1519;
  wire T1520;
  wire T1521;
  wire T1522;
  wire T1523;
  wire T1524;
  wire T1525;
  wire T1526;
  wire T1527;
  wire T1528;
  wire T1529;
  wire T1530;
  wire T1531;
  wire T1532;
  wire T1533;
  wire T1534;
  wire T1535;
  wire T1536;
  wire T1537;
  wire T1538;
  wire T1539;
  wire[54:0] T3174;
  wire[30:0] T1540;
  wire[30:0] T1541;
  wire[8:0] T1542;
  wire[4:0] T1543;
  wire[3:0] T1544;
  wire[21:0] T1545;
  wire[4:0] T1546;
  wire[16:0] T1547;
  wire T1548;
  wire T1549;
  wire T1550;
  wire T1551;
  wire flitsAreTail_1;
  wire T1552;
  wire T1553;
  wire T1554;
  wire T1555;
  wire[53:0] T1556;
  wire T1557;
  wire[30:0] T1558;
  wire T1559;
  wire T1560;
  wire T1561;
  wire T1562;
  wire T1563;
  wire[54:0] T1564;
  wire[54:0] T1565;
  wire T1566;
  wire T1567;
  wire T1568;
  wire T1569;
  wire T1570;
  wire T1571;
  wire T1572;
  wire T1573;
  wire T1574;
  wire T1575;
  wire[54:0] T1576;
  wire[54:0] T1577;
  wire T3175;
  reg [54:0] R1578;
  wire[54:0] T3176;
  wire[54:0] T1579;
  wire[54:0] T3177;
  wire T1580;
  wire T1581;
  wire[54:0] T1582;
  wire[54:0] T1583;
  wire T1584;
  wire T1585;
  wire[1:0] T1586;
  wire[1:0] T1587;
  wire[1:0] T1588;
  wire T1589;
  wire[2:0] T1590;
  reg [2:0] R1591;
  wire[2:0] T3178;
  wire[1:0] T1592;
  wire T1593;
  wire T1594;
  wire T1595;
  wire T1596;
  wire T1597;
  wire T1598;
  wire T1599;
  wire T1600;
  wire T1601;
  wire[2:0] T1602;
  wire T1603;
  wire T1604;
  wire T1605;
  wire T1606;
  wire T1607;
  wire T1608;
  wire T1609;
  wire T1610;
  wire T1611;
  wire T1612;
  wire T1613;
  wire T1614;
  wire T1615;
  wire T3179;
  wire T1616;
  wire T1617;
  wire[3:0] T1618;
  wire[3:0] T1619;
  wire[3:0] T1620;
  wire T1621;
  wire[2:0] T1622;
  wire[3:0] T1623;
  wire T1624;
  wire T1625;
  wire T1626;
  wire T1627;
  wire T1628;
  wire T1629;
  wire T1630;
  wire[2:0] T1631;
  wire T1632;
  wire T1633;
  wire T1634;
  wire T1635;
  wire T1636;
  wire T1637;
  wire T1638;
  wire T1639;
  wire[53:0] T1640;
  wire T1641;
  wire[30:0] T1642;
  wire T1643;
  wire T1644;
  reg  R1645;
  wire T3180;
  wire[2:0] T1646;
  wire[30:0] T1647;
  wire[54:0] T1648;
  wire[1:0] T1649;
  wire[1:0] T1650;
  wire[1:0] T1651;
  wire[3:0] T1652;
  wire T1653;
  wire T1654;
  wire[15:0] T1655;
  wire T1656;
  wire T1657;
  wire T1658;
  wire T1659;
  wire T1660;
  wire T1661;
  wire T1662;
  wire T1663;
  wire T1664;
  wire T1665;
  wire T1666;
  wire T1667;
  wire T1668;
  wire T1669;
  wire T1670;
  wire T1671;
  wire T1672;
  wire T1673;
  wire T1674;
  wire T1675;
  wire T1676;
  wire T1677;
  wire T1678;
  wire T1679;
  wire T1680;
  wire T1681;
  wire T1682;
  wire T1683;
  wire[54:0] T3181;
  wire[30:0] T1684;
  wire[30:0] T1685;
  wire[8:0] T1686;
  wire[4:0] T1687;
  wire[3:0] T1688;
  wire[21:0] T1689;
  wire[4:0] T1690;
  wire[16:0] T1691;
  wire T1692;
  wire T1693;
  wire T1694;
  wire T1695;
  wire flitsAreTail_0;
  wire T1696;
  wire T1697;
  wire T1698;
  wire T1699;
  wire[53:0] T1700;
  wire T1701;
  wire[30:0] T1702;
  wire T1703;
  wire T1704;
  wire T1705;
  wire T1706;
  wire T1707;
  wire[54:0] T1708;
  wire[54:0] T1709;
  wire T1710;
  wire T1711;
  wire T1712;
  wire T1713;
  wire T1714;
  wire T1715;
  wire T1716;
  wire T1717;
  wire T1718;
  wire T1719;
  wire T1720;
  wire T1721;
  wire T1722;
  wire[9:0] T1723;
  wire[9:0] T1724;
  wire[4:0] T1725;
  wire[2:0] T1726;
  wire[1:0] T1727;
  wire readyToXmit_0_4;
  wire T1728;
  wire T1729;
  wire T1730;
  wire T1731;
  wire T1732;
  wire T1733;
  wire T1734;
  wire T1735;
  wire[7:0] T1736;
  wire[2:0] T1737;
  wire T1738;
  wire T1739;
  wire T1740;
  wire T1741;
  wire T1742;
  wire T1743;
  wire T1744;
  wire readyToXmit_1_4;
  wire T1745;
  wire T1746;
  wire T1747;
  wire T1748;
  wire T1749;
  wire T1750;
  wire T1751;
  wire T1752;
  wire[7:0] T1753;
  wire[2:0] T1754;
  wire T1755;
  wire T1756;
  wire T1757;
  wire T1758;
  wire T1759;
  wire T1760;
  wire T1761;
  wire readyToXmit_2_4;
  wire T1762;
  wire T1763;
  wire T1764;
  wire T1765;
  wire T1766;
  wire T1767;
  wire T1768;
  wire T1769;
  wire[7:0] T1770;
  wire[2:0] T1771;
  wire T1772;
  wire T1773;
  wire T1774;
  wire T1775;
  wire T1776;
  wire T1777;
  wire T1778;
  wire[1:0] T1779;
  wire readyToXmit_3_4;
  wire T1780;
  wire T1781;
  wire T1782;
  wire T1783;
  wire T1784;
  wire T1785;
  wire T1786;
  wire T1787;
  wire[7:0] T1788;
  wire[2:0] T1789;
  wire T1790;
  wire T1791;
  wire T1792;
  wire T1793;
  wire T1794;
  wire T1795;
  wire T1796;
  wire readyToXmit_4_4;
  wire T1797;
  wire T1798;
  wire T1799;
  wire T1800;
  wire T1801;
  wire T1802;
  wire T1803;
  wire T1804;
  wire[7:0] T1805;
  wire[2:0] T1806;
  wire T1807;
  wire T1808;
  wire T1809;
  wire T1810;
  wire T1811;
  wire T1812;
  wire T1813;
  wire[4:0] T1814;
  wire[2:0] T1815;
  wire[1:0] T1816;
  wire readyToXmit_5_4;
  wire T1817;
  wire T1818;
  wire T1819;
  wire T1820;
  wire T1821;
  wire T1822;
  wire T1823;
  wire T1824;
  wire[7:0] T1825;
  wire[2:0] T1826;
  wire T1827;
  wire T1828;
  wire T1829;
  wire T1830;
  wire T1831;
  wire T1832;
  wire T1833;
  wire readyToXmit_6_4;
  wire T1834;
  wire T1835;
  wire T1836;
  wire T1837;
  wire T1838;
  wire T1839;
  wire T1840;
  wire T1841;
  wire[7:0] T1842;
  wire[2:0] T1843;
  wire T1844;
  wire T1845;
  wire T1846;
  wire T1847;
  wire T1848;
  wire T1849;
  wire T1850;
  wire readyToXmit_7_4;
  wire T1851;
  wire T1852;
  wire T1853;
  wire T1854;
  wire T1855;
  wire T1856;
  wire T1857;
  wire T1858;
  wire[7:0] T1859;
  wire[2:0] T1860;
  wire T1861;
  wire T1862;
  wire T1863;
  wire T1864;
  wire T1865;
  wire T1866;
  wire T1867;
  wire[1:0] T1868;
  wire readyToXmit_8_4;
  wire T1869;
  wire T1870;
  wire T1871;
  wire T1872;
  wire T1873;
  wire T1874;
  wire T1875;
  wire T1876;
  wire[7:0] T1877;
  wire[2:0] T1878;
  wire T1879;
  wire T1880;
  wire T1881;
  wire T1882;
  wire T1883;
  wire T1884;
  wire T1885;
  wire readyToXmit_9_4;
  wire T1886;
  wire T1887;
  wire T1888;
  wire T1889;
  wire T1890;
  wire T1891;
  wire T1892;
  wire T1893;
  wire[7:0] T1894;
  wire[2:0] T1895;
  wire T1896;
  wire T1897;
  wire T1898;
  wire T1899;
  wire T1900;
  wire T1901;
  wire T1902;
  wire T1903;
  wire T1904;
  wire T1905;
  wire[9:0] T1906;
  wire[9:0] T1907;
  wire[4:0] T1908;
  wire[2:0] T1909;
  wire[1:0] T1910;
  wire readyToXmit_0_3;
  wire T1911;
  wire T1912;
  wire T1913;
  wire T1914;
  wire T1915;
  wire readyToXmit_1_3;
  wire T1916;
  wire T1917;
  wire T1918;
  wire T1919;
  wire T1920;
  wire readyToXmit_2_3;
  wire T1921;
  wire T1922;
  wire T1923;
  wire T1924;
  wire T1925;
  wire[1:0] T1926;
  wire readyToXmit_3_3;
  wire T1927;
  wire T1928;
  wire T1929;
  wire T1930;
  wire T1931;
  wire readyToXmit_4_3;
  wire T1932;
  wire T1933;
  wire T1934;
  wire T1935;
  wire T1936;
  wire[4:0] T1937;
  wire[2:0] T1938;
  wire[1:0] T1939;
  wire readyToXmit_5_3;
  wire T1940;
  wire T1941;
  wire T1942;
  wire T1943;
  wire T1944;
  wire readyToXmit_6_3;
  wire T1945;
  wire T1946;
  wire T1947;
  wire T1948;
  wire T1949;
  wire readyToXmit_7_3;
  wire T1950;
  wire T1951;
  wire T1952;
  wire T1953;
  wire T1954;
  wire[1:0] T1955;
  wire readyToXmit_8_3;
  wire T1956;
  wire T1957;
  wire T1958;
  wire T1959;
  wire T1960;
  wire readyToXmit_9_3;
  wire T1961;
  wire T1962;
  wire T1963;
  wire T1964;
  wire T1965;
  wire T1966;
  wire T1967;
  wire T1968;
  wire[9:0] T1969;
  wire[9:0] T1970;
  wire[4:0] T1971;
  wire[2:0] T1972;
  wire[1:0] T1973;
  wire readyToXmit_0_2;
  wire T1974;
  wire T1975;
  wire T1976;
  wire T1977;
  wire T1978;
  wire readyToXmit_1_2;
  wire T1979;
  wire T1980;
  wire T1981;
  wire T1982;
  wire T1983;
  wire readyToXmit_2_2;
  wire T1984;
  wire T1985;
  wire T1986;
  wire T1987;
  wire T1988;
  wire[1:0] T1989;
  wire readyToXmit_3_2;
  wire T1990;
  wire T1991;
  wire T1992;
  wire T1993;
  wire T1994;
  wire readyToXmit_4_2;
  wire T1995;
  wire T1996;
  wire T1997;
  wire T1998;
  wire T1999;
  wire[4:0] T2000;
  wire[2:0] T2001;
  wire[1:0] T2002;
  wire readyToXmit_5_2;
  wire T2003;
  wire T2004;
  wire T2005;
  wire T2006;
  wire T2007;
  wire readyToXmit_6_2;
  wire T2008;
  wire T2009;
  wire T2010;
  wire T2011;
  wire T2012;
  wire readyToXmit_7_2;
  wire T2013;
  wire T2014;
  wire T2015;
  wire T2016;
  wire T2017;
  wire[1:0] T2018;
  wire readyToXmit_8_2;
  wire T2019;
  wire T2020;
  wire T2021;
  wire T2022;
  wire T2023;
  wire readyToXmit_9_2;
  wire T2024;
  wire T2025;
  wire T2026;
  wire T2027;
  wire T2028;
  wire T2029;
  wire T2030;
  wire T2031;
  wire[9:0] T2032;
  wire[9:0] T2033;
  wire[4:0] T2034;
  wire[2:0] T2035;
  wire[1:0] T2036;
  wire readyToXmit_0_1;
  wire T2037;
  wire T2038;
  wire T2039;
  wire T2040;
  wire T2041;
  wire readyToXmit_1_1;
  wire T2042;
  wire T2043;
  wire T2044;
  wire T2045;
  wire T2046;
  wire readyToXmit_2_1;
  wire T2047;
  wire T2048;
  wire T2049;
  wire T2050;
  wire T2051;
  wire[1:0] T2052;
  wire readyToXmit_3_1;
  wire T2053;
  wire T2054;
  wire T2055;
  wire T2056;
  wire T2057;
  wire readyToXmit_4_1;
  wire T2058;
  wire T2059;
  wire T2060;
  wire T2061;
  wire T2062;
  wire[4:0] T2063;
  wire[2:0] T2064;
  wire[1:0] T2065;
  wire readyToXmit_5_1;
  wire T2066;
  wire T2067;
  wire T2068;
  wire T2069;
  wire T2070;
  wire readyToXmit_6_1;
  wire T2071;
  wire T2072;
  wire T2073;
  wire T2074;
  wire T2075;
  wire readyToXmit_7_1;
  wire T2076;
  wire T2077;
  wire T2078;
  wire T2079;
  wire T2080;
  wire[1:0] T2081;
  wire readyToXmit_8_1;
  wire T2082;
  wire T2083;
  wire T2084;
  wire T2085;
  wire T2086;
  wire readyToXmit_9_1;
  wire T2087;
  wire T2088;
  wire T2089;
  wire T2090;
  wire T2091;
  wire T2092;
  wire T2093;
  wire T2094;
  wire[9:0] T2095;
  wire[9:0] T2096;
  wire[4:0] T2097;
  wire[2:0] T2098;
  wire[1:0] T2099;
  wire readyToXmit_0_0;
  wire T2100;
  wire T2101;
  wire T2102;
  wire T2103;
  wire T2104;
  wire readyToXmit_1_0;
  wire T2105;
  wire T2106;
  wire T2107;
  wire T2108;
  wire T2109;
  wire readyToXmit_2_0;
  wire T2110;
  wire T2111;
  wire T2112;
  wire T2113;
  wire T2114;
  wire[1:0] T2115;
  wire readyToXmit_3_0;
  wire T2116;
  wire T2117;
  wire T2118;
  wire T2119;
  wire T2120;
  wire readyToXmit_4_0;
  wire T2121;
  wire T2122;
  wire T2123;
  wire T2124;
  wire T2125;
  wire[4:0] T2126;
  wire[2:0] T2127;
  wire[1:0] T2128;
  wire readyToXmit_5_0;
  wire T2129;
  wire T2130;
  wire T2131;
  wire T2132;
  wire T2133;
  wire readyToXmit_6_0;
  wire T2134;
  wire T2135;
  wire T2136;
  wire T2137;
  wire T2138;
  wire readyToXmit_7_0;
  wire T2139;
  wire T2140;
  wire T2141;
  wire T2142;
  wire T2143;
  wire[1:0] T2144;
  wire readyToXmit_8_0;
  wire T2145;
  wire T2146;
  wire T2147;
  wire T2148;
  wire T2149;
  wire readyToXmit_9_0;
  wire T2150;
  wire T2151;
  wire T2152;
  wire T2153;
  wire T2154;
  wire T2155;
  wire T2156;
  wire T2157;
  wire T2158;
  wire T2159;
  wire T2160;
  wire T2161;
  wire T2162;
  wire T2163;
  wire T2164;
  wire T2165;
  wire T2166;
  wire T2167;
  wire T2168;
  wire T2169;
  wire T2170;
  wire T2171;
  wire T2172;
  wire T2173;
  wire T2174;
  wire T2175;
  reg [1:0] validVCs_0_0;
  reg  R2176;
  wire T2177;
  wire T2178;
  wire T2179;
  wire T2180;
  reg  R2181;
  wire T2182;
  wire T2183;
  wire T2184;
  wire T2185;
  reg [1:0] validVCs_0_1;
  reg  R2186;
  wire T2187;
  wire T2188;
  wire T2189;
  wire T2190;
  reg  R2191;
  wire T2192;
  wire T2193;
  wire T2194;
  wire T2195;
  reg [1:0] validVCs_0_2;
  reg  R2196;
  wire T2197;
  wire T2198;
  wire T2199;
  wire T2200;
  reg  R2201;
  wire T2202;
  wire T2203;
  wire T2204;
  wire T2205;
  reg [1:0] validVCs_0_3;
  reg  R2206;
  wire T2207;
  wire T2208;
  wire T2209;
  wire T2210;
  reg  R2211;
  wire T2212;
  wire T2213;
  wire T2214;
  wire T2215;
  reg [1:0] validVCs_0_4;
  reg  R2216;
  wire T2217;
  wire T2218;
  wire T2219;
  wire T2220;
  reg  R2221;
  wire T2222;
  wire T2223;
  wire T2224;
  wire T2225;
  reg [1:0] validVCs_1_0;
  reg  R2226;
  wire T2227;
  wire T2228;
  wire T2229;
  wire T2230;
  reg  R2231;
  wire T2232;
  wire T2233;
  wire T2234;
  wire T2235;
  reg [1:0] validVCs_1_1;
  reg  R2236;
  wire T2237;
  wire T2238;
  wire T2239;
  wire T2240;
  reg  R2241;
  wire T2242;
  wire T2243;
  wire T2244;
  wire T2245;
  reg [1:0] validVCs_1_2;
  reg  R2246;
  wire T2247;
  wire T2248;
  wire T2249;
  wire T2250;
  reg  R2251;
  wire T2252;
  wire T2253;
  wire T2254;
  wire T2255;
  reg [1:0] validVCs_1_3;
  reg  R2256;
  wire T2257;
  wire T2258;
  wire T2259;
  wire T2260;
  reg  R2261;
  wire T2262;
  wire T2263;
  wire T2264;
  wire T2265;
  reg [1:0] validVCs_1_4;
  reg  R2266;
  wire T2267;
  wire T2268;
  wire T2269;
  wire T2270;
  reg  R2271;
  wire T2272;
  wire T2273;
  wire T2274;
  wire T2275;
  reg [1:0] validVCs_2_0;
  reg  R2276;
  wire T2277;
  wire T2278;
  wire T2279;
  wire T2280;
  reg  R2281;
  wire T2282;
  wire T2283;
  wire T2284;
  wire T2285;
  reg [1:0] validVCs_2_1;
  reg  R2286;
  wire T2287;
  wire T2288;
  wire T2289;
  wire T2290;
  reg  R2291;
  wire T2292;
  wire T2293;
  wire T2294;
  wire T2295;
  reg [1:0] validVCs_2_2;
  reg  R2296;
  wire T2297;
  wire T2298;
  wire T2299;
  wire T2300;
  reg  R2301;
  wire T2302;
  wire T2303;
  wire T2304;
  wire T2305;
  reg [1:0] validVCs_2_3;
  reg  R2306;
  wire T2307;
  wire T2308;
  wire T2309;
  wire T2310;
  reg  R2311;
  wire T2312;
  wire T2313;
  wire T2314;
  wire T2315;
  reg [1:0] validVCs_2_4;
  reg  R2316;
  wire T2317;
  wire T2318;
  wire T2319;
  wire T2320;
  reg  R2321;
  wire T2322;
  wire T2323;
  wire T2324;
  wire T2325;
  reg [1:0] validVCs_3_0;
  reg  R2326;
  wire T2327;
  wire T2328;
  wire T2329;
  wire T2330;
  reg  R2331;
  wire T2332;
  wire T2333;
  wire T2334;
  wire T2335;
  reg [1:0] validVCs_3_1;
  reg  R2336;
  wire T2337;
  wire T2338;
  wire T2339;
  wire T2340;
  reg  R2341;
  wire T2342;
  wire T2343;
  wire T2344;
  wire T2345;
  reg [1:0] validVCs_3_2;
  reg  R2346;
  wire T2347;
  wire T2348;
  wire T2349;
  wire T2350;
  reg  R2351;
  wire T2352;
  wire T2353;
  wire T2354;
  wire T2355;
  reg [1:0] validVCs_3_3;
  reg  R2356;
  wire T2357;
  wire T2358;
  wire T2359;
  wire T2360;
  reg  R2361;
  wire T2362;
  wire T2363;
  wire T2364;
  wire T2365;
  reg [1:0] validVCs_3_4;
  reg  R2366;
  wire T2367;
  wire T2368;
  wire T2369;
  wire T2370;
  reg  R2371;
  wire T2372;
  wire T2373;
  wire T2374;
  wire T2375;
  reg [1:0] validVCs_4_0;
  reg  R2376;
  wire T2377;
  wire T2378;
  wire T2379;
  wire T2380;
  reg  R2381;
  wire T2382;
  wire T2383;
  wire T2384;
  wire T2385;
  reg [1:0] validVCs_4_1;
  reg  R2386;
  wire T2387;
  wire T2388;
  wire T2389;
  wire T2390;
  reg  R2391;
  wire T2392;
  wire T2393;
  wire T2394;
  wire T2395;
  reg [1:0] validVCs_4_2;
  reg  R2396;
  wire T2397;
  wire T2398;
  wire T2399;
  wire T2400;
  reg  R2401;
  wire T2402;
  wire T2403;
  wire T2404;
  wire T2405;
  reg [1:0] validVCs_4_3;
  reg  R2406;
  wire T2407;
  wire T2408;
  wire T2409;
  wire T2410;
  reg  R2411;
  wire T2412;
  wire T2413;
  wire T2414;
  wire T2415;
  reg [1:0] validVCs_4_4;
  reg  R2416;
  wire T2417;
  wire T2418;
  wire T2419;
  wire T2420;
  reg  R2421;
  wire T2422;
  wire T2423;
  wire T2424;
  wire T2425;
  reg [1:0] validVCs_5_0;
  reg  R2426;
  wire T2427;
  wire T2428;
  wire T2429;
  wire T2430;
  reg  R2431;
  wire T2432;
  wire T2433;
  wire T2434;
  wire T2435;
  reg [1:0] validVCs_5_1;
  reg  R2436;
  wire T2437;
  wire T2438;
  wire T2439;
  wire T2440;
  reg  R2441;
  wire T2442;
  wire T2443;
  wire T2444;
  wire T2445;
  reg [1:0] validVCs_5_2;
  reg  R2446;
  wire T2447;
  wire T2448;
  wire T2449;
  wire T2450;
  reg  R2451;
  wire T2452;
  wire T2453;
  wire T2454;
  wire T2455;
  reg [1:0] validVCs_5_3;
  reg  R2456;
  wire T2457;
  wire T2458;
  wire T2459;
  wire T2460;
  reg  R2461;
  wire T2462;
  wire T2463;
  wire T2464;
  wire T2465;
  reg [1:0] validVCs_5_4;
  reg  R2466;
  wire T2467;
  wire T2468;
  wire T2469;
  wire T2470;
  reg  R2471;
  wire T2472;
  wire T2473;
  wire T2474;
  wire T2475;
  reg [1:0] validVCs_6_0;
  reg  R2476;
  wire T2477;
  wire T2478;
  wire T2479;
  wire T2480;
  reg  R2481;
  wire T2482;
  wire T2483;
  wire T2484;
  wire T2485;
  reg [1:0] validVCs_6_1;
  reg  R2486;
  wire T2487;
  wire T2488;
  wire T2489;
  wire T2490;
  reg  R2491;
  wire T2492;
  wire T2493;
  wire T2494;
  wire T2495;
  reg [1:0] validVCs_6_2;
  reg  R2496;
  wire T2497;
  wire T2498;
  wire T2499;
  wire T2500;
  reg  R2501;
  wire T2502;
  wire T2503;
  wire T2504;
  wire T2505;
  reg [1:0] validVCs_6_3;
  reg  R2506;
  wire T2507;
  wire T2508;
  wire T2509;
  wire T2510;
  reg  R2511;
  wire T2512;
  wire T2513;
  wire T2514;
  wire T2515;
  reg [1:0] validVCs_6_4;
  reg  R2516;
  wire T2517;
  wire T2518;
  wire T2519;
  wire T2520;
  reg  R2521;
  wire T2522;
  wire T2523;
  wire T2524;
  wire T2525;
  reg [1:0] validVCs_7_0;
  reg  R2526;
  wire T2527;
  wire T2528;
  wire T2529;
  wire T2530;
  reg  R2531;
  wire T2532;
  wire T2533;
  wire T2534;
  wire T2535;
  reg [1:0] validVCs_7_1;
  reg  R2536;
  wire T2537;
  wire T2538;
  wire T2539;
  wire T2540;
  reg  R2541;
  wire T2542;
  wire T2543;
  wire T2544;
  wire T2545;
  reg [1:0] validVCs_7_2;
  reg  R2546;
  wire T2547;
  wire T2548;
  wire T2549;
  wire T2550;
  reg  R2551;
  wire T2552;
  wire T2553;
  wire T2554;
  wire T2555;
  reg [1:0] validVCs_7_3;
  reg  R2556;
  wire T2557;
  wire T2558;
  wire T2559;
  wire T2560;
  reg  R2561;
  wire T2562;
  wire T2563;
  wire T2564;
  wire T2565;
  reg [1:0] validVCs_7_4;
  reg  R2566;
  wire T2567;
  wire T2568;
  wire T2569;
  wire T2570;
  reg  R2571;
  wire T2572;
  wire T2573;
  wire T2574;
  wire T2575;
  reg [1:0] validVCs_8_0;
  reg  R2576;
  wire T2577;
  wire T2578;
  wire T2579;
  wire T2580;
  reg  R2581;
  wire T2582;
  wire T2583;
  wire T2584;
  wire T2585;
  reg [1:0] validVCs_8_1;
  reg  R2586;
  wire T2587;
  wire T2588;
  wire T2589;
  wire T2590;
  reg  R2591;
  wire T2592;
  wire T2593;
  wire T2594;
  wire T2595;
  reg [1:0] validVCs_8_2;
  reg  R2596;
  wire T2597;
  wire T2598;
  wire T2599;
  wire T2600;
  reg  R2601;
  wire T2602;
  wire T2603;
  wire T2604;
  wire T2605;
  reg [1:0] validVCs_8_3;
  reg  R2606;
  wire T2607;
  wire T2608;
  wire T2609;
  wire T2610;
  reg  R2611;
  wire T2612;
  wire T2613;
  wire T2614;
  wire T2615;
  reg [1:0] validVCs_8_4;
  reg  R2616;
  wire T2617;
  wire T2618;
  wire T2619;
  wire T2620;
  reg  R2621;
  wire T2622;
  wire T2623;
  wire T2624;
  wire T2625;
  reg [1:0] validVCs_9_0;
  reg  R2626;
  wire T2627;
  wire T2628;
  wire T2629;
  wire T2630;
  reg  R2631;
  wire T2632;
  wire T2633;
  wire T2634;
  wire T2635;
  reg [1:0] validVCs_9_1;
  reg  R2636;
  wire T2637;
  wire T2638;
  wire T2639;
  wire T2640;
  reg  R2641;
  wire T2642;
  wire T2643;
  wire T2644;
  wire T2645;
  reg [1:0] validVCs_9_2;
  reg  R2646;
  wire T2647;
  wire T2648;
  wire T2649;
  wire T2650;
  reg  R2651;
  wire T2652;
  wire T2653;
  wire T2654;
  wire T2655;
  reg [1:0] validVCs_9_3;
  reg  R2656;
  wire T2657;
  wire T2658;
  wire T2659;
  wire T2660;
  reg  R2661;
  wire T2662;
  wire T2663;
  wire T2664;
  wire T2665;
  reg [1:0] validVCs_9_4;
  reg  R2666;
  wire T2667;
  wire T2668;
  wire T2669;
  wire T2670;
  reg  R2671;
  wire T2672;
  wire T2673;
  wire T2674;
  reg [2:0] R2675;
  wire[2:0] T3182;
  wire[2:0] T2676;
  wire[2:0] T2677;
  wire[30:0] T2678;
  wire T2679;
  wire T2680;
  wire T2681;
  wire T2682;
  reg [7:0] R2683;
  wire[7:0] T3183;
  wire[7:0] T2684;
  wire T2685;
  wire T2686;
  wire T2687;
  reg  R2688;
  wire T3184;
  reg [2:0] R2689;
  wire[2:0] T3185;
  wire[2:0] T2690;
  wire[2:0] T2691;
  wire[30:0] T2692;
  wire T2693;
  wire T2694;
  wire T2695;
  wire T2696;
  reg [7:0] R2697;
  wire[7:0] T3186;
  wire[7:0] T2698;
  wire T2699;
  wire T2700;
  wire T2701;
  reg  R2702;
  wire T3187;
  reg [2:0] R2703;
  wire[2:0] T3188;
  wire[2:0] T2704;
  wire[2:0] T2705;
  wire[30:0] T2706;
  wire T2707;
  wire T2708;
  wire T2709;
  wire T2710;
  reg [7:0] R2711;
  wire[7:0] T3189;
  wire[7:0] T2712;
  wire T2713;
  wire T2714;
  wire T2715;
  reg  R2716;
  wire T3190;
  reg [2:0] R2717;
  wire[2:0] T3191;
  wire[2:0] T2718;
  wire[2:0] T2719;
  wire[30:0] T2720;
  wire T2721;
  wire T2722;
  wire T2723;
  wire T2724;
  reg [7:0] R2725;
  wire[7:0] T3192;
  wire[7:0] T2726;
  wire T2727;
  wire T2728;
  wire T2729;
  reg  R2730;
  wire T3193;
  reg [2:0] R2731;
  wire[2:0] T3194;
  wire[2:0] T2732;
  wire[2:0] T2733;
  wire[30:0] T2734;
  wire T2735;
  wire T2736;
  wire T2737;
  wire T2738;
  reg [7:0] R2739;
  wire[7:0] T3195;
  wire[7:0] T2740;
  wire T2741;
  wire T2742;
  wire T2743;
  reg  R2744;
  wire T3196;
  reg [2:0] R2745;
  wire[2:0] T3197;
  wire[2:0] T2746;
  wire[2:0] T2747;
  wire[30:0] T2748;
  wire T2749;
  wire T2750;
  wire T2751;
  wire T2752;
  reg [7:0] R2753;
  wire[7:0] T3198;
  wire[7:0] T2754;
  wire T2755;
  wire T2756;
  wire T2757;
  reg  R2758;
  wire T3199;
  reg [2:0] R2759;
  wire[2:0] T3200;
  wire[2:0] T2760;
  wire[2:0] T2761;
  wire[30:0] T2762;
  wire T2763;
  wire T2764;
  wire T2765;
  wire T2766;
  reg [7:0] R2767;
  wire[7:0] T3201;
  wire[7:0] T2768;
  wire T2769;
  wire T2770;
  wire T2771;
  reg  R2772;
  wire T3202;
  reg [2:0] R2773;
  wire[2:0] T3203;
  wire[2:0] T2774;
  wire[2:0] T2775;
  wire[30:0] T2776;
  wire T2777;
  wire T2778;
  wire T2779;
  wire T2780;
  reg [7:0] R2781;
  wire[7:0] T3204;
  wire[7:0] T2782;
  wire T2783;
  wire T2784;
  wire T2785;
  reg  R2786;
  wire T3205;
  reg [2:0] R2787;
  wire[2:0] T3206;
  wire[2:0] T2788;
  wire[2:0] T2789;
  wire[30:0] T2790;
  wire T2791;
  wire T2792;
  wire T2793;
  wire T2794;
  reg [7:0] R2795;
  wire[7:0] T3207;
  wire[7:0] T2796;
  wire T2797;
  wire T2798;
  wire T2799;
  reg  R2800;
  wire T3208;
  reg [2:0] R2801;
  wire[2:0] T3209;
  wire[2:0] T2802;
  wire[2:0] T2803;
  wire[30:0] T2804;
  wire T2805;
  wire T2806;
  wire T2807;
  wire T2808;
  reg [7:0] R2809;
  wire[7:0] T3210;
  wire[7:0] T2810;
  wire T2811;
  wire T2812;
  wire T2813;
  reg  R2814;
  wire T3211;
  wire T2815;
  wire T2816;
  wire T2817;
  wire T2818;
  wire T2819;
  wire T2820;
  wire T2821;
  wire T2822;
  wire T2823;
  wire T2824;
  wire T2825;
  wire T2826;
  wire T2827;
  wire T2828;
  wire T2829;
  wire T2830;
  wire T2831;
  wire T2832;
  wire T2833;
  wire T2834;
  wire T2835;
  wire T2836;
  wire T2837;
  wire T2838;
  wire T2839;
  wire T2840;
  wire T2841;
  wire T2842;
  wire T2843;
  wire T2844;
  wire T2845;
  wire T2846;
  wire T2847;
  wire T2848;
  wire T2849;
  wire T2850;
  wire T2851;
  wire T2852;
  wire T2853;
  wire T2854;
  wire T2855;
  wire T2856;
  wire T2857;
  wire T2858;
  wire T2859;
  wire T2860;
  wire T2861;
  wire T2862;
  wire T2863;
  wire T2864;
  wire T2865;
  wire T2866;
  wire T2867;
  wire T2868;
  wire T2869;
  wire T2870;
  wire T2871;
  wire T2872;
  wire T2873;
  wire T2874;
  wire T2875;
  wire T2876;
  wire T2877;
  wire T2878;
  wire T2879;
  wire T2880;
  wire T2881;
  wire T2882;
  wire T2883;
  wire T2884;
  wire T2885;
  wire T2886;
  wire T2887;
  wire T2888;
  wire T2889;
  wire T2890;
  wire T2891;
  wire T2892;
  wire T2893;
  wire T2894;
  wire T2895;
  wire T2896;
  wire T2897;
  wire T2898;
  wire T2899;
  wire T2900;
  wire T2901;
  wire T2902;
  wire T2903;
  wire T2904;
  wire T2905;
  wire T2906;
  wire T2907;
  wire T2908;
  wire T2909;
  wire T2910;
  wire T2911;
  wire T2912;
  wire T2913;
  wire T2914;
  wire T2915;
  wire T2916;
  wire T2917;
  wire T2918;
  wire T2919;
  wire T2920;
  wire T2921;
  wire T2922;
  wire T2923;
  wire T2924;
  wire T2925;
  wire T2926;
  wire T2927;
  wire T2928;
  wire T2929;
  wire T2930;
  wire T2931;
  wire T2932;
  wire T2933;
  wire T2934;
  wire T2935;
  wire T2936;
  wire T2937;
  wire T2938;
  wire T2939;
  wire T2940;
  wire T2941;
  wire T2942;
  wire T2943;
  wire T2944;
  wire T2945;
  wire T2946;
  wire T2947;
  wire T2948;
  wire T2949;
  wire T2950;
  wire T2951;
  wire T2952;
  wire T2953;
  wire T2954;
  wire T2955;
  wire T2956;
  wire T2957;
  wire T2958;
  wire T2959;
  wire T2960;
  wire T2961;
  wire T2962;
  wire T2963;
  wire T2964;
  wire T2965;
  wire T2966;
  wire T2967;
  wire T2968;
  wire T2969;
  wire T2970;
  wire T2971;
  wire T2972;
  wire T2973;
  wire T2974;
  wire T2975;
  wire T2976;
  wire T2977;
  wire T2978;
  wire T2979;
  wire T2980;
  wire T2981;
  wire T2982;
  wire T2983;
  wire T2984;
  wire T2985;
  wire T2986;
  wire T2987;
  wire T2988;
  wire T2989;
  wire T2990;
  wire T2991;
  wire T2992;
  wire T2993;
  wire T2994;
  wire T2995;
  wire T2996;
  wire T2997;
  wire T2998;
  wire T2999;
  wire T3000;
  wire T3001;
  wire T3002;
  wire T3003;
  wire T3004;
  wire T3005;
  wire T3006;
  wire T3007;
  wire T3008;
  wire T3009;
  wire T3010;
  wire T3011;
  wire T3012;
  wire T3013;
  wire T3014;
  wire T3015;
  wire T3016;
  wire T3017;
  wire T3018;
  wire T3019;
  wire T3020;
  wire T3021;
  wire T3022;
  wire T3023;
  wire T3024;
  wire T3025;
  wire T3026;
  wire T3027;
  wire T3028;
  wire T3029;
  wire T3030;
  wire T3031;
  wire T3032;
  wire T3033;
  wire T3034;
  wire T3035;
  wire T3036;
  wire T3037;
  wire T3038;
  wire T3039;
  wire T3040;
  wire T3041;
  wire T3042;
  wire T3043;
  wire T3044;
  wire T3045;
  wire T3046;
  wire T3047;
  wire T3048;
  wire T3049;
  wire T3050;
  wire T3051;
  wire T3052;
  wire T3053;
  wire T3054;
  wire T3055;
  wire T3056;
  wire T3057;
  wire T3058;
  wire T3059;
  wire T3060;
  wire T3061;
  wire T3062;
  wire T3063;
  wire T3064;
  wire T3065;
  wire T3066;
  wire T3067;
  wire T3068;
  wire T3069;
  wire T3070;
  wire T3071;
  wire T3072;
  wire T3073;
  wire T3074;
  wire T3075;
  wire T3076;
  wire T3077;
  wire T3078;
  wire T3079;
  wire T3080;
  wire T3081;
  wire T3082;
  wire T3083;
  wire T3084;
  wire T3085;
  wire T3086;
  wire T3087;
  wire T3088;
  wire T3089;
  wire T3090;
  wire T3091;
  wire T3092;
  wire T3093;
  wire T3094;
  wire[31:0] T3212;
  wire T3095;
  wire T3096;
  reg  R3097;
  reg [54:0] R3098;
  wire[54:0] T3099;
  wire[54:0] T3213;
  reg  R3100;
  reg [54:0] R3101;
  wire[54:0] T3102;
  wire[54:0] T3214;
  reg  R3103;
  reg [54:0] R3104;
  wire[54:0] T3105;
  wire[54:0] T3215;
  reg  R3106;
  reg [54:0] R3107;
  wire[54:0] T3108;
  wire[54:0] T3216;
  reg  R3109;
  reg [54:0] R3110;
  wire[54:0] T3111;
  wire[54:0] T3217;
  wire[1:0] VCRouterOutputStateManagement_io_currentState;
  wire[1:0] VCRouterOutputStateManagement_1_io_currentState;
  wire[1:0] VCRouterOutputStateManagement_2_io_currentState;
  wire[1:0] VCRouterOutputStateManagement_3_io_currentState;
  wire[1:0] VCRouterOutputStateManagement_4_io_currentState;
  wire CreditGen_io_outCredit_grant;
  wire[54:0] RouterRegFile_io_readData;
  wire RouterRegFile_io_readValid;
  wire[54:0] RouterRegFile_io_readPipelineReg_1;
  wire[54:0] RouterRegFile_io_readPipelineReg_0;
  wire RouterRegFile_io_rvPipelineReg_1;
  wire RouterRegFile_io_rvPipelineReg_0;
  wire[15:0] CMeshDOR_io_outHeadFlit_packetID;
  wire CMeshDOR_io_outHeadFlit_isTail;
  wire CMeshDOR_io_outHeadFlit_vcPort;
  wire[3:0] CMeshDOR_io_outHeadFlit_packetType;
  wire[1:0] CMeshDOR_io_outHeadFlit_destination_2;
  wire[1:0] CMeshDOR_io_outHeadFlit_destination_1;
  wire[1:0] CMeshDOR_io_outHeadFlit_destination_0;
  wire[2:0] CMeshDOR_io_outHeadFlit_priorityLevel;
  wire[2:0] CMeshDOR_io_result;
  wire[1:0] CMeshDOR_io_vcsAvailable_4;
  wire[1:0] CMeshDOR_io_vcsAvailable_3;
  wire[1:0] CMeshDOR_io_vcsAvailable_2;
  wire[1:0] CMeshDOR_io_vcsAvailable_1;
  wire[1:0] CMeshDOR_io_vcsAvailable_0;
  wire[2:0] VCRouterStateManagement_io_currentState;
  wire CreditGen_1_io_outCredit_grant;
  wire[54:0] RouterRegFile_1_io_readData;
  wire RouterRegFile_1_io_readValid;
  wire[54:0] RouterRegFile_1_io_readPipelineReg_1;
  wire[54:0] RouterRegFile_1_io_readPipelineReg_0;
  wire RouterRegFile_1_io_rvPipelineReg_1;
  wire RouterRegFile_1_io_rvPipelineReg_0;
  wire[15:0] CMeshDOR_1_io_outHeadFlit_packetID;
  wire CMeshDOR_1_io_outHeadFlit_isTail;
  wire CMeshDOR_1_io_outHeadFlit_vcPort;
  wire[3:0] CMeshDOR_1_io_outHeadFlit_packetType;
  wire[1:0] CMeshDOR_1_io_outHeadFlit_destination_2;
  wire[1:0] CMeshDOR_1_io_outHeadFlit_destination_1;
  wire[1:0] CMeshDOR_1_io_outHeadFlit_destination_0;
  wire[2:0] CMeshDOR_1_io_outHeadFlit_priorityLevel;
  wire[2:0] CMeshDOR_1_io_result;
  wire[1:0] CMeshDOR_1_io_vcsAvailable_4;
  wire[1:0] CMeshDOR_1_io_vcsAvailable_3;
  wire[1:0] CMeshDOR_1_io_vcsAvailable_2;
  wire[1:0] CMeshDOR_1_io_vcsAvailable_1;
  wire[1:0] CMeshDOR_1_io_vcsAvailable_0;
  wire[2:0] VCRouterStateManagement_1_io_currentState;
  wire CreditGen_2_io_outCredit_grant;
  wire[54:0] RouterRegFile_2_io_readData;
  wire RouterRegFile_2_io_readValid;
  wire[54:0] RouterRegFile_2_io_readPipelineReg_1;
  wire[54:0] RouterRegFile_2_io_readPipelineReg_0;
  wire RouterRegFile_2_io_rvPipelineReg_1;
  wire RouterRegFile_2_io_rvPipelineReg_0;
  wire[15:0] CMeshDOR_2_io_outHeadFlit_packetID;
  wire CMeshDOR_2_io_outHeadFlit_isTail;
  wire CMeshDOR_2_io_outHeadFlit_vcPort;
  wire[3:0] CMeshDOR_2_io_outHeadFlit_packetType;
  wire[1:0] CMeshDOR_2_io_outHeadFlit_destination_2;
  wire[1:0] CMeshDOR_2_io_outHeadFlit_destination_1;
  wire[1:0] CMeshDOR_2_io_outHeadFlit_destination_0;
  wire[2:0] CMeshDOR_2_io_outHeadFlit_priorityLevel;
  wire[2:0] CMeshDOR_2_io_result;
  wire[1:0] CMeshDOR_2_io_vcsAvailable_4;
  wire[1:0] CMeshDOR_2_io_vcsAvailable_3;
  wire[1:0] CMeshDOR_2_io_vcsAvailable_2;
  wire[1:0] CMeshDOR_2_io_vcsAvailable_1;
  wire[1:0] CMeshDOR_2_io_vcsAvailable_0;
  wire[2:0] VCRouterStateManagement_2_io_currentState;
  wire CreditGen_3_io_outCredit_grant;
  wire[54:0] RouterRegFile_3_io_readData;
  wire RouterRegFile_3_io_readValid;
  wire[54:0] RouterRegFile_3_io_readPipelineReg_1;
  wire[54:0] RouterRegFile_3_io_readPipelineReg_0;
  wire RouterRegFile_3_io_rvPipelineReg_1;
  wire RouterRegFile_3_io_rvPipelineReg_0;
  wire[15:0] CMeshDOR_3_io_outHeadFlit_packetID;
  wire CMeshDOR_3_io_outHeadFlit_isTail;
  wire CMeshDOR_3_io_outHeadFlit_vcPort;
  wire[3:0] CMeshDOR_3_io_outHeadFlit_packetType;
  wire[1:0] CMeshDOR_3_io_outHeadFlit_destination_2;
  wire[1:0] CMeshDOR_3_io_outHeadFlit_destination_1;
  wire[1:0] CMeshDOR_3_io_outHeadFlit_destination_0;
  wire[2:0] CMeshDOR_3_io_outHeadFlit_priorityLevel;
  wire[2:0] CMeshDOR_3_io_result;
  wire[1:0] CMeshDOR_3_io_vcsAvailable_4;
  wire[1:0] CMeshDOR_3_io_vcsAvailable_3;
  wire[1:0] CMeshDOR_3_io_vcsAvailable_2;
  wire[1:0] CMeshDOR_3_io_vcsAvailable_1;
  wire[1:0] CMeshDOR_3_io_vcsAvailable_0;
  wire[2:0] VCRouterStateManagement_3_io_currentState;
  wire CreditGen_4_io_outCredit_grant;
  wire[54:0] RouterRegFile_4_io_readData;
  wire RouterRegFile_4_io_readValid;
  wire[54:0] RouterRegFile_4_io_readPipelineReg_1;
  wire[54:0] RouterRegFile_4_io_readPipelineReg_0;
  wire RouterRegFile_4_io_rvPipelineReg_1;
  wire RouterRegFile_4_io_rvPipelineReg_0;
  wire[15:0] CMeshDOR_4_io_outHeadFlit_packetID;
  wire CMeshDOR_4_io_outHeadFlit_isTail;
  wire CMeshDOR_4_io_outHeadFlit_vcPort;
  wire[3:0] CMeshDOR_4_io_outHeadFlit_packetType;
  wire[1:0] CMeshDOR_4_io_outHeadFlit_destination_2;
  wire[1:0] CMeshDOR_4_io_outHeadFlit_destination_1;
  wire[1:0] CMeshDOR_4_io_outHeadFlit_destination_0;
  wire[2:0] CMeshDOR_4_io_outHeadFlit_priorityLevel;
  wire[2:0] CMeshDOR_4_io_result;
  wire[1:0] CMeshDOR_4_io_vcsAvailable_4;
  wire[1:0] CMeshDOR_4_io_vcsAvailable_3;
  wire[1:0] CMeshDOR_4_io_vcsAvailable_2;
  wire[1:0] CMeshDOR_4_io_vcsAvailable_1;
  wire[1:0] CMeshDOR_4_io_vcsAvailable_0;
  wire[2:0] VCRouterStateManagement_4_io_currentState;
  wire CreditGen_5_io_outCredit_grant;
  wire[54:0] RouterRegFile_5_io_readData;
  wire RouterRegFile_5_io_readValid;
  wire[54:0] RouterRegFile_5_io_readPipelineReg_1;
  wire[54:0] RouterRegFile_5_io_readPipelineReg_0;
  wire RouterRegFile_5_io_rvPipelineReg_1;
  wire RouterRegFile_5_io_rvPipelineReg_0;
  wire[15:0] CMeshDOR_5_io_outHeadFlit_packetID;
  wire CMeshDOR_5_io_outHeadFlit_isTail;
  wire CMeshDOR_5_io_outHeadFlit_vcPort;
  wire[3:0] CMeshDOR_5_io_outHeadFlit_packetType;
  wire[1:0] CMeshDOR_5_io_outHeadFlit_destination_2;
  wire[1:0] CMeshDOR_5_io_outHeadFlit_destination_1;
  wire[1:0] CMeshDOR_5_io_outHeadFlit_destination_0;
  wire[2:0] CMeshDOR_5_io_outHeadFlit_priorityLevel;
  wire[2:0] CMeshDOR_5_io_result;
  wire[1:0] CMeshDOR_5_io_vcsAvailable_4;
  wire[1:0] CMeshDOR_5_io_vcsAvailable_3;
  wire[1:0] CMeshDOR_5_io_vcsAvailable_2;
  wire[1:0] CMeshDOR_5_io_vcsAvailable_1;
  wire[1:0] CMeshDOR_5_io_vcsAvailable_0;
  wire[2:0] VCRouterStateManagement_5_io_currentState;
  wire CreditGen_6_io_outCredit_grant;
  wire[54:0] RouterRegFile_6_io_readData;
  wire RouterRegFile_6_io_readValid;
  wire[54:0] RouterRegFile_6_io_readPipelineReg_1;
  wire[54:0] RouterRegFile_6_io_readPipelineReg_0;
  wire RouterRegFile_6_io_rvPipelineReg_1;
  wire RouterRegFile_6_io_rvPipelineReg_0;
  wire[15:0] CMeshDOR_6_io_outHeadFlit_packetID;
  wire CMeshDOR_6_io_outHeadFlit_isTail;
  wire CMeshDOR_6_io_outHeadFlit_vcPort;
  wire[3:0] CMeshDOR_6_io_outHeadFlit_packetType;
  wire[1:0] CMeshDOR_6_io_outHeadFlit_destination_2;
  wire[1:0] CMeshDOR_6_io_outHeadFlit_destination_1;
  wire[1:0] CMeshDOR_6_io_outHeadFlit_destination_0;
  wire[2:0] CMeshDOR_6_io_outHeadFlit_priorityLevel;
  wire[2:0] CMeshDOR_6_io_result;
  wire[1:0] CMeshDOR_6_io_vcsAvailable_4;
  wire[1:0] CMeshDOR_6_io_vcsAvailable_3;
  wire[1:0] CMeshDOR_6_io_vcsAvailable_2;
  wire[1:0] CMeshDOR_6_io_vcsAvailable_1;
  wire[1:0] CMeshDOR_6_io_vcsAvailable_0;
  wire[2:0] VCRouterStateManagement_6_io_currentState;
  wire CreditGen_7_io_outCredit_grant;
  wire[54:0] RouterRegFile_7_io_readData;
  wire RouterRegFile_7_io_readValid;
  wire[54:0] RouterRegFile_7_io_readPipelineReg_1;
  wire[54:0] RouterRegFile_7_io_readPipelineReg_0;
  wire RouterRegFile_7_io_rvPipelineReg_1;
  wire RouterRegFile_7_io_rvPipelineReg_0;
  wire[15:0] CMeshDOR_7_io_outHeadFlit_packetID;
  wire CMeshDOR_7_io_outHeadFlit_isTail;
  wire CMeshDOR_7_io_outHeadFlit_vcPort;
  wire[3:0] CMeshDOR_7_io_outHeadFlit_packetType;
  wire[1:0] CMeshDOR_7_io_outHeadFlit_destination_2;
  wire[1:0] CMeshDOR_7_io_outHeadFlit_destination_1;
  wire[1:0] CMeshDOR_7_io_outHeadFlit_destination_0;
  wire[2:0] CMeshDOR_7_io_outHeadFlit_priorityLevel;
  wire[2:0] CMeshDOR_7_io_result;
  wire[1:0] CMeshDOR_7_io_vcsAvailable_4;
  wire[1:0] CMeshDOR_7_io_vcsAvailable_3;
  wire[1:0] CMeshDOR_7_io_vcsAvailable_2;
  wire[1:0] CMeshDOR_7_io_vcsAvailable_1;
  wire[1:0] CMeshDOR_7_io_vcsAvailable_0;
  wire[2:0] VCRouterStateManagement_7_io_currentState;
  wire CreditGen_8_io_outCredit_grant;
  wire[54:0] RouterRegFile_8_io_readData;
  wire RouterRegFile_8_io_readValid;
  wire[54:0] RouterRegFile_8_io_readPipelineReg_1;
  wire[54:0] RouterRegFile_8_io_readPipelineReg_0;
  wire RouterRegFile_8_io_rvPipelineReg_1;
  wire RouterRegFile_8_io_rvPipelineReg_0;
  wire[15:0] CMeshDOR_8_io_outHeadFlit_packetID;
  wire CMeshDOR_8_io_outHeadFlit_isTail;
  wire CMeshDOR_8_io_outHeadFlit_vcPort;
  wire[3:0] CMeshDOR_8_io_outHeadFlit_packetType;
  wire[1:0] CMeshDOR_8_io_outHeadFlit_destination_2;
  wire[1:0] CMeshDOR_8_io_outHeadFlit_destination_1;
  wire[1:0] CMeshDOR_8_io_outHeadFlit_destination_0;
  wire[2:0] CMeshDOR_8_io_outHeadFlit_priorityLevel;
  wire[2:0] CMeshDOR_8_io_result;
  wire[1:0] CMeshDOR_8_io_vcsAvailable_4;
  wire[1:0] CMeshDOR_8_io_vcsAvailable_3;
  wire[1:0] CMeshDOR_8_io_vcsAvailable_2;
  wire[1:0] CMeshDOR_8_io_vcsAvailable_1;
  wire[1:0] CMeshDOR_8_io_vcsAvailable_0;
  wire[2:0] VCRouterStateManagement_8_io_currentState;
  wire CreditGen_9_io_outCredit_grant;
  wire[54:0] RouterRegFile_9_io_readData;
  wire RouterRegFile_9_io_readValid;
  wire[54:0] RouterRegFile_9_io_readPipelineReg_1;
  wire[54:0] RouterRegFile_9_io_readPipelineReg_0;
  wire RouterRegFile_9_io_rvPipelineReg_1;
  wire RouterRegFile_9_io_rvPipelineReg_0;
  wire[15:0] CMeshDOR_9_io_outHeadFlit_packetID;
  wire CMeshDOR_9_io_outHeadFlit_isTail;
  wire CMeshDOR_9_io_outHeadFlit_vcPort;
  wire[3:0] CMeshDOR_9_io_outHeadFlit_packetType;
  wire[1:0] CMeshDOR_9_io_outHeadFlit_destination_2;
  wire[1:0] CMeshDOR_9_io_outHeadFlit_destination_1;
  wire[1:0] CMeshDOR_9_io_outHeadFlit_destination_0;
  wire[2:0] CMeshDOR_9_io_outHeadFlit_priorityLevel;
  wire[2:0] CMeshDOR_9_io_result;
  wire[1:0] CMeshDOR_9_io_vcsAvailable_4;
  wire[1:0] CMeshDOR_9_io_vcsAvailable_3;
  wire[1:0] CMeshDOR_9_io_vcsAvailable_2;
  wire[1:0] CMeshDOR_9_io_vcsAvailable_1;
  wire[1:0] CMeshDOR_9_io_vcsAvailable_0;
  wire[2:0] VCRouterStateManagement_9_io_currentState;
  wire CreditCon_io_outCredit;
  wire CreditCon_1_io_outCredit;
  wire CreditCon_2_io_outCredit;
  wire CreditCon_3_io_outCredit;
  wire CreditCon_4_io_outCredit;
  wire CreditCon_5_io_outCredit;
  wire CreditCon_6_io_outCredit;
  wire CreditCon_7_io_outCredit;
  wire CreditCon_8_io_outCredit;
  wire CreditCon_9_io_outCredit;
  wire[54:0] switch_io_outPorts_4_x;
  wire[54:0] switch_io_outPorts_3_x;
  wire[54:0] switch_io_outPorts_2_x;
  wire[54:0] switch_io_outPorts_1_x;
  wire[54:0] switch_io_outPorts_0_x;
  wire swAllocator_io_requests_4_9_grant;
  wire swAllocator_io_requests_4_8_grant;
  wire swAllocator_io_requests_4_7_grant;
  wire swAllocator_io_requests_4_6_grant;
  wire swAllocator_io_requests_4_5_grant;
  wire swAllocator_io_requests_4_4_grant;
  wire swAllocator_io_requests_4_3_grant;
  wire swAllocator_io_requests_4_2_grant;
  wire swAllocator_io_requests_4_1_grant;
  wire swAllocator_io_requests_4_0_grant;
  wire swAllocator_io_requests_3_9_grant;
  wire swAllocator_io_requests_3_8_grant;
  wire swAllocator_io_requests_3_7_grant;
  wire swAllocator_io_requests_3_6_grant;
  wire swAllocator_io_requests_3_5_grant;
  wire swAllocator_io_requests_3_4_grant;
  wire swAllocator_io_requests_3_3_grant;
  wire swAllocator_io_requests_3_2_grant;
  wire swAllocator_io_requests_3_1_grant;
  wire swAllocator_io_requests_3_0_grant;
  wire swAllocator_io_requests_2_9_grant;
  wire swAllocator_io_requests_2_8_grant;
  wire swAllocator_io_requests_2_7_grant;
  wire swAllocator_io_requests_2_6_grant;
  wire swAllocator_io_requests_2_5_grant;
  wire swAllocator_io_requests_2_4_grant;
  wire swAllocator_io_requests_2_3_grant;
  wire swAllocator_io_requests_2_2_grant;
  wire swAllocator_io_requests_2_1_grant;
  wire swAllocator_io_requests_2_0_grant;
  wire swAllocator_io_requests_1_9_grant;
  wire swAllocator_io_requests_1_8_grant;
  wire swAllocator_io_requests_1_7_grant;
  wire swAllocator_io_requests_1_6_grant;
  wire swAllocator_io_requests_1_5_grant;
  wire swAllocator_io_requests_1_4_grant;
  wire swAllocator_io_requests_1_3_grant;
  wire swAllocator_io_requests_1_2_grant;
  wire swAllocator_io_requests_1_1_grant;
  wire swAllocator_io_requests_1_0_grant;
  wire swAllocator_io_requests_0_9_grant;
  wire swAllocator_io_requests_0_8_grant;
  wire swAllocator_io_requests_0_7_grant;
  wire swAllocator_io_requests_0_6_grant;
  wire swAllocator_io_requests_0_5_grant;
  wire swAllocator_io_requests_0_4_grant;
  wire swAllocator_io_requests_0_3_grant;
  wire swAllocator_io_requests_0_2_grant;
  wire swAllocator_io_requests_0_1_grant;
  wire swAllocator_io_requests_0_0_grant;
  wire[3:0] swAllocator_io_chosens_4;
  wire[3:0] swAllocator_io_chosens_3;
  wire[3:0] swAllocator_io_chosens_2;
  wire[3:0] swAllocator_io_chosens_1;
  wire[3:0] swAllocator_io_chosens_0;
  wire vcAllocator_io_resources_9_valid;
  wire vcAllocator_io_resources_8_valid;
  wire vcAllocator_io_resources_7_valid;
  wire vcAllocator_io_resources_6_valid;
  wire vcAllocator_io_resources_5_valid;
  wire vcAllocator_io_resources_4_valid;
  wire vcAllocator_io_resources_3_valid;
  wire vcAllocator_io_resources_2_valid;
  wire vcAllocator_io_resources_1_valid;
  wire vcAllocator_io_resources_0_valid;
  wire[3:0] vcAllocator_io_chosens_9;
  wire[3:0] vcAllocator_io_chosens_8;
  wire[3:0] vcAllocator_io_chosens_7;
  wire[3:0] vcAllocator_io_chosens_6;
  wire[3:0] vcAllocator_io_chosens_5;
  wire[3:0] vcAllocator_io_chosens_4;
  wire[3:0] vcAllocator_io_chosens_3;
  wire[3:0] vcAllocator_io_chosens_2;
  wire[3:0] vcAllocator_io_chosens_1;
  wire[3:0] vcAllocator_io_chosens_0;
  wire RouterBuffer_io_enq_ready;
  wire RouterBuffer_io_deq_valid;
  wire[54:0] RouterBuffer_io_deq_bits_x;
  wire[54:0] ReplaceVCPort_io_newFlit_x;
  wire RouterBuffer_1_io_enq_ready;
  wire RouterBuffer_1_io_deq_valid;
  wire[54:0] RouterBuffer_1_io_deq_bits_x;
  wire[54:0] ReplaceVCPort_1_io_newFlit_x;
  wire RouterBuffer_2_io_enq_ready;
  wire RouterBuffer_2_io_deq_valid;
  wire[54:0] RouterBuffer_2_io_deq_bits_x;
  wire[54:0] ReplaceVCPort_2_io_newFlit_x;
  wire RouterBuffer_3_io_enq_ready;
  wire RouterBuffer_3_io_deq_valid;
  wire[54:0] RouterBuffer_3_io_deq_bits_x;
  wire[54:0] ReplaceVCPort_3_io_newFlit_x;
  wire RouterBuffer_4_io_enq_ready;
  wire RouterBuffer_4_io_deq_valid;
  wire[54:0] RouterBuffer_4_io_deq_bits_x;
  wire[54:0] ReplaceVCPort_4_io_newFlit_x;
  wire RouterBuffer_5_io_enq_ready;
  wire RouterBuffer_5_io_deq_valid;
  wire[54:0] RouterBuffer_5_io_deq_bits_x;
  wire[54:0] ReplaceVCPort_5_io_newFlit_x;
  wire RouterBuffer_6_io_enq_ready;
  wire RouterBuffer_6_io_deq_valid;
  wire[54:0] RouterBuffer_6_io_deq_bits_x;
  wire[54:0] ReplaceVCPort_6_io_newFlit_x;
  wire RouterBuffer_7_io_enq_ready;
  wire RouterBuffer_7_io_deq_valid;
  wire[54:0] RouterBuffer_7_io_deq_bits_x;
  wire[54:0] ReplaceVCPort_7_io_newFlit_x;
  wire RouterBuffer_8_io_enq_ready;
  wire RouterBuffer_8_io_deq_valid;
  wire[54:0] RouterBuffer_8_io_deq_bits_x;
  wire[54:0] ReplaceVCPort_8_io_newFlit_x;
  wire RouterBuffer_9_io_enq_ready;
  wire RouterBuffer_9_io_deq_valid;
  wire[54:0] RouterBuffer_9_io_deq_bits_x;
  wire[54:0] ReplaceVCPort_9_io_newFlit_x;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    T0 = 1'b0;
    T17 = 1'b0;
    T22 = 1'b0;
    T39 = 1'b0;
    T44 = 1'b0;
    T61 = 1'b0;
    T66 = 1'b0;
    T83 = 1'b0;
    T88 = 1'b0;
    T105 = 1'b0;
    T110 = 1'b0;
    T127 = 1'b0;
    T132 = 1'b0;
    T149 = 1'b0;
    T154 = 1'b0;
    T171 = 1'b0;
    T176 = 1'b0;
    T193 = 1'b0;
    T198 = 1'b0;
    T215 = 1'b0;
    R282 = {2{1'b0}};
    R295 = {1{1'b0}};
    R349 = {1{1'b0}};
    R426 = {2{1'b0}};
    R439 = {1{1'b0}};
    R493 = {1{1'b0}};
    R570 = {2{1'b0}};
    R583 = {1{1'b0}};
    R637 = {1{1'b0}};
    R714 = {2{1'b0}};
    R727 = {1{1'b0}};
    R781 = {1{1'b0}};
    R858 = {2{1'b0}};
    R871 = {1{1'b0}};
    R925 = {1{1'b0}};
    R1002 = {2{1'b0}};
    R1015 = {1{1'b0}};
    R1069 = {1{1'b0}};
    R1146 = {2{1'b0}};
    R1159 = {1{1'b0}};
    R1213 = {1{1'b0}};
    R1290 = {2{1'b0}};
    R1303 = {1{1'b0}};
    R1357 = {1{1'b0}};
    R1434 = {2{1'b0}};
    R1447 = {1{1'b0}};
    R1501 = {1{1'b0}};
    R1578 = {2{1'b0}};
    R1591 = {1{1'b0}};
    R1645 = {1{1'b0}};
    validVCs_0_0 = {1{1'b0}};
    R2176 = {1{1'b0}};
    R2181 = {1{1'b0}};
    validVCs_0_1 = {1{1'b0}};
    R2186 = {1{1'b0}};
    R2191 = {1{1'b0}};
    validVCs_0_2 = {1{1'b0}};
    R2196 = {1{1'b0}};
    R2201 = {1{1'b0}};
    validVCs_0_3 = {1{1'b0}};
    R2206 = {1{1'b0}};
    R2211 = {1{1'b0}};
    validVCs_0_4 = {1{1'b0}};
    R2216 = {1{1'b0}};
    R2221 = {1{1'b0}};
    validVCs_1_0 = {1{1'b0}};
    R2226 = {1{1'b0}};
    R2231 = {1{1'b0}};
    validVCs_1_1 = {1{1'b0}};
    R2236 = {1{1'b0}};
    R2241 = {1{1'b0}};
    validVCs_1_2 = {1{1'b0}};
    R2246 = {1{1'b0}};
    R2251 = {1{1'b0}};
    validVCs_1_3 = {1{1'b0}};
    R2256 = {1{1'b0}};
    R2261 = {1{1'b0}};
    validVCs_1_4 = {1{1'b0}};
    R2266 = {1{1'b0}};
    R2271 = {1{1'b0}};
    validVCs_2_0 = {1{1'b0}};
    R2276 = {1{1'b0}};
    R2281 = {1{1'b0}};
    validVCs_2_1 = {1{1'b0}};
    R2286 = {1{1'b0}};
    R2291 = {1{1'b0}};
    validVCs_2_2 = {1{1'b0}};
    R2296 = {1{1'b0}};
    R2301 = {1{1'b0}};
    validVCs_2_3 = {1{1'b0}};
    R2306 = {1{1'b0}};
    R2311 = {1{1'b0}};
    validVCs_2_4 = {1{1'b0}};
    R2316 = {1{1'b0}};
    R2321 = {1{1'b0}};
    validVCs_3_0 = {1{1'b0}};
    R2326 = {1{1'b0}};
    R2331 = {1{1'b0}};
    validVCs_3_1 = {1{1'b0}};
    R2336 = {1{1'b0}};
    R2341 = {1{1'b0}};
    validVCs_3_2 = {1{1'b0}};
    R2346 = {1{1'b0}};
    R2351 = {1{1'b0}};
    validVCs_3_3 = {1{1'b0}};
    R2356 = {1{1'b0}};
    R2361 = {1{1'b0}};
    validVCs_3_4 = {1{1'b0}};
    R2366 = {1{1'b0}};
    R2371 = {1{1'b0}};
    validVCs_4_0 = {1{1'b0}};
    R2376 = {1{1'b0}};
    R2381 = {1{1'b0}};
    validVCs_4_1 = {1{1'b0}};
    R2386 = {1{1'b0}};
    R2391 = {1{1'b0}};
    validVCs_4_2 = {1{1'b0}};
    R2396 = {1{1'b0}};
    R2401 = {1{1'b0}};
    validVCs_4_3 = {1{1'b0}};
    R2406 = {1{1'b0}};
    R2411 = {1{1'b0}};
    validVCs_4_4 = {1{1'b0}};
    R2416 = {1{1'b0}};
    R2421 = {1{1'b0}};
    validVCs_5_0 = {1{1'b0}};
    R2426 = {1{1'b0}};
    R2431 = {1{1'b0}};
    validVCs_5_1 = {1{1'b0}};
    R2436 = {1{1'b0}};
    R2441 = {1{1'b0}};
    validVCs_5_2 = {1{1'b0}};
    R2446 = {1{1'b0}};
    R2451 = {1{1'b0}};
    validVCs_5_3 = {1{1'b0}};
    R2456 = {1{1'b0}};
    R2461 = {1{1'b0}};
    validVCs_5_4 = {1{1'b0}};
    R2466 = {1{1'b0}};
    R2471 = {1{1'b0}};
    validVCs_6_0 = {1{1'b0}};
    R2476 = {1{1'b0}};
    R2481 = {1{1'b0}};
    validVCs_6_1 = {1{1'b0}};
    R2486 = {1{1'b0}};
    R2491 = {1{1'b0}};
    validVCs_6_2 = {1{1'b0}};
    R2496 = {1{1'b0}};
    R2501 = {1{1'b0}};
    validVCs_6_3 = {1{1'b0}};
    R2506 = {1{1'b0}};
    R2511 = {1{1'b0}};
    validVCs_6_4 = {1{1'b0}};
    R2516 = {1{1'b0}};
    R2521 = {1{1'b0}};
    validVCs_7_0 = {1{1'b0}};
    R2526 = {1{1'b0}};
    R2531 = {1{1'b0}};
    validVCs_7_1 = {1{1'b0}};
    R2536 = {1{1'b0}};
    R2541 = {1{1'b0}};
    validVCs_7_2 = {1{1'b0}};
    R2546 = {1{1'b0}};
    R2551 = {1{1'b0}};
    validVCs_7_3 = {1{1'b0}};
    R2556 = {1{1'b0}};
    R2561 = {1{1'b0}};
    validVCs_7_4 = {1{1'b0}};
    R2566 = {1{1'b0}};
    R2571 = {1{1'b0}};
    validVCs_8_0 = {1{1'b0}};
    R2576 = {1{1'b0}};
    R2581 = {1{1'b0}};
    validVCs_8_1 = {1{1'b0}};
    R2586 = {1{1'b0}};
    R2591 = {1{1'b0}};
    validVCs_8_2 = {1{1'b0}};
    R2596 = {1{1'b0}};
    R2601 = {1{1'b0}};
    validVCs_8_3 = {1{1'b0}};
    R2606 = {1{1'b0}};
    R2611 = {1{1'b0}};
    validVCs_8_4 = {1{1'b0}};
    R2616 = {1{1'b0}};
    R2621 = {1{1'b0}};
    validVCs_9_0 = {1{1'b0}};
    R2626 = {1{1'b0}};
    R2631 = {1{1'b0}};
    validVCs_9_1 = {1{1'b0}};
    R2636 = {1{1'b0}};
    R2641 = {1{1'b0}};
    validVCs_9_2 = {1{1'b0}};
    R2646 = {1{1'b0}};
    R2651 = {1{1'b0}};
    validVCs_9_3 = {1{1'b0}};
    R2656 = {1{1'b0}};
    R2661 = {1{1'b0}};
    validVCs_9_4 = {1{1'b0}};
    R2666 = {1{1'b0}};
    R2671 = {1{1'b0}};
    R2675 = {1{1'b0}};
    R2683 = {1{1'b0}};
    R2688 = {1{1'b0}};
    R2689 = {1{1'b0}};
    R2697 = {1{1'b0}};
    R2702 = {1{1'b0}};
    R2703 = {1{1'b0}};
    R2711 = {1{1'b0}};
    R2716 = {1{1'b0}};
    R2717 = {1{1'b0}};
    R2725 = {1{1'b0}};
    R2730 = {1{1'b0}};
    R2731 = {1{1'b0}};
    R2739 = {1{1'b0}};
    R2744 = {1{1'b0}};
    R2745 = {1{1'b0}};
    R2753 = {1{1'b0}};
    R2758 = {1{1'b0}};
    R2759 = {1{1'b0}};
    R2767 = {1{1'b0}};
    R2772 = {1{1'b0}};
    R2773 = {1{1'b0}};
    R2781 = {1{1'b0}};
    R2786 = {1{1'b0}};
    R2787 = {1{1'b0}};
    R2795 = {1{1'b0}};
    R2800 = {1{1'b0}};
    R2801 = {1{1'b0}};
    R2809 = {1{1'b0}};
    R2814 = {1{1'b0}};
    R3097 = {1{1'b0}};
    R3098 = {2{1'b0}};
    R3100 = {1{1'b0}};
    R3101 = {2{1'b0}};
    R3103 = {1{1'b0}};
    R3104 = {2{1'b0}};
    R3106 = {1{1'b0}};
    R3107 = {2{1'b0}};
    R3109 = {1{1'b0}};
    R3110 = {2{1'b0}};
  end
// synthesis translate_on
`endif

`ifndef SYNTHESIS
// synthesis translate_off
//  assign io_counters_0_counterIndex = {1{1'b0}};
//  assign io_counters_1_counterIndex = {1{1'b0}};
//  assign io_counters_1_counterVal = {1{1'b0}};
// synthesis translate_on
`endif
  assign T1 = T2 | reset;
  assign T2 = T13 | T3;
  assign T3 = ~ T4;
  assign T4 = T5 == 1'h1;
  assign T5 = T6;
  assign T6 = T11 ? T9 : T7;
  assign T7 = T8[6'h24:6'h24];
  assign T8 = io_inChannels_4_flit_x[6'h36:1'h1];
  assign T9 = T10[4'hd:4'hd];
  assign T10 = io_inChannels_4_flit_x[5'h1f:1'h1];
  assign T11 = T12 == 1'h1;
  assign T12 = io_inChannels_4_flit_x[1'h0:1'h0];
  assign T13 = T15 | T14;
  assign T14 = ~ io_inChannels_4_flitValid;
  assign T15 = T16 & T4;
  assign T16 = RouterBuffer_9_io_enq_ready & io_inChannels_4_flitValid;
  assign T18 = T19 | reset;
  assign T19 = T21 | T20;
  assign T20 = T379 & T4;
  assign T21 = ~ T379;
  assign T23 = T24 | reset;
  assign T24 = T35 | T25;
  assign T25 = ~ T26;
  assign T26 = T27 == 1'h0;
  assign T27 = T28;
  assign T28 = T33 ? T31 : T29;
  assign T29 = T30[6'h24:6'h24];
  assign T30 = io_inChannels_4_flit_x[6'h36:1'h1];
  assign T31 = T32[4'hd:4'hd];
  assign T32 = io_inChannels_4_flit_x[5'h1f:1'h1];
  assign T33 = T34 == 1'h1;
  assign T34 = io_inChannels_4_flit_x[1'h0:1'h0];
  assign T35 = T37 | T36;
  assign T36 = ~ io_inChannels_4_flitValid;
  assign T37 = T38 & T26;
  assign T38 = RouterBuffer_8_io_enq_ready & io_inChannels_4_flitValid;
  assign T40 = T41 | reset;
  assign T41 = T43 | T42;
  assign T42 = T523 & T26;
  assign T43 = ~ T523;
  assign T45 = T46 | reset;
  assign T46 = T57 | T47;
  assign T47 = ~ T48;
  assign T48 = T49 == 1'h1;
  assign T49 = T50;
  assign T50 = T55 ? T53 : T51;
  assign T51 = T52[6'h24:6'h24];
  assign T52 = io_inChannels_3_flit_x[6'h36:1'h1];
  assign T53 = T54[4'hd:4'hd];
  assign T54 = io_inChannels_3_flit_x[5'h1f:1'h1];
  assign T55 = T56 == 1'h1;
  assign T56 = io_inChannels_3_flit_x[1'h0:1'h0];
  assign T57 = T59 | T58;
  assign T58 = ~ io_inChannels_3_flitValid;
  assign T59 = T60 & T48;
  assign T60 = RouterBuffer_7_io_enq_ready & io_inChannels_3_flitValid;
  assign T62 = T63 | reset;
  assign T63 = T65 | T64;
  assign T64 = T667 & T48;
  assign T65 = ~ T667;
  assign T67 = T68 | reset;
  assign T68 = T79 | T69;
  assign T69 = ~ T70;
  assign T70 = T71 == 1'h0;
  assign T71 = T72;
  assign T72 = T77 ? T75 : T73;
  assign T73 = T74[6'h24:6'h24];
  assign T74 = io_inChannels_3_flit_x[6'h36:1'h1];
  assign T75 = T76[4'hd:4'hd];
  assign T76 = io_inChannels_3_flit_x[5'h1f:1'h1];
  assign T77 = T78 == 1'h1;
  assign T78 = io_inChannels_3_flit_x[1'h0:1'h0];
  assign T79 = T81 | T80;
  assign T80 = ~ io_inChannels_3_flitValid;
  assign T81 = T82 & T70;
  assign T82 = RouterBuffer_6_io_enq_ready & io_inChannels_3_flitValid;
  assign T84 = T85 | reset;
  assign T85 = T87 | T86;
  assign T86 = T811 & T70;
  assign T87 = ~ T811;
  assign T89 = T90 | reset;
  assign T90 = T101 | T91;
  assign T91 = ~ T92;
  assign T92 = T93 == 1'h1;
  assign T93 = T94;
  assign T94 = T99 ? T97 : T95;
  assign T95 = T96[6'h24:6'h24];
  assign T96 = io_inChannels_2_flit_x[6'h36:1'h1];
  assign T97 = T98[4'hd:4'hd];
  assign T98 = io_inChannels_2_flit_x[5'h1f:1'h1];
  assign T99 = T100 == 1'h1;
  assign T100 = io_inChannels_2_flit_x[1'h0:1'h0];
  assign T101 = T103 | T102;
  assign T102 = ~ io_inChannels_2_flitValid;
  assign T103 = T104 & T92;
  assign T104 = RouterBuffer_5_io_enq_ready & io_inChannels_2_flitValid;
  assign T106 = T107 | reset;
  assign T107 = T109 | T108;
  assign T108 = T955 & T92;
  assign T109 = ~ T955;
  assign T111 = T112 | reset;
  assign T112 = T123 | T113;
  assign T113 = ~ T114;
  assign T114 = T115 == 1'h0;
  assign T115 = T116;
  assign T116 = T121 ? T119 : T117;
  assign T117 = T118[6'h24:6'h24];
  assign T118 = io_inChannels_2_flit_x[6'h36:1'h1];
  assign T119 = T120[4'hd:4'hd];
  assign T120 = io_inChannels_2_flit_x[5'h1f:1'h1];
  assign T121 = T122 == 1'h1;
  assign T122 = io_inChannels_2_flit_x[1'h0:1'h0];
  assign T123 = T125 | T124;
  assign T124 = ~ io_inChannels_2_flitValid;
  assign T125 = T126 & T114;
  assign T126 = RouterBuffer_4_io_enq_ready & io_inChannels_2_flitValid;
  assign T128 = T129 | reset;
  assign T129 = T131 | T130;
  assign T130 = T1099 & T114;
  assign T131 = ~ T1099;
  assign T133 = T134 | reset;
  assign T134 = T145 | T135;
  assign T135 = ~ T136;
  assign T136 = T137 == 1'h1;
  assign T137 = T138;
  assign T138 = T143 ? T141 : T139;
  assign T139 = T140[6'h24:6'h24];
  assign T140 = io_inChannels_1_flit_x[6'h36:1'h1];
  assign T141 = T142[4'hd:4'hd];
  assign T142 = io_inChannels_1_flit_x[5'h1f:1'h1];
  assign T143 = T144 == 1'h1;
  assign T144 = io_inChannels_1_flit_x[1'h0:1'h0];
  assign T145 = T147 | T146;
  assign T146 = ~ io_inChannels_1_flitValid;
  assign T147 = T148 & T136;
  assign T148 = RouterBuffer_3_io_enq_ready & io_inChannels_1_flitValid;
  assign T150 = T151 | reset;
  assign T151 = T153 | T152;
  assign T152 = T1243 & T136;
  assign T153 = ~ T1243;
  assign T155 = T156 | reset;
  assign T156 = T167 | T157;
  assign T157 = ~ T158;
  assign T158 = T159 == 1'h0;
  assign T159 = T160;
  assign T160 = T165 ? T163 : T161;
  assign T161 = T162[6'h24:6'h24];
  assign T162 = io_inChannels_1_flit_x[6'h36:1'h1];
  assign T163 = T164[4'hd:4'hd];
  assign T164 = io_inChannels_1_flit_x[5'h1f:1'h1];
  assign T165 = T166 == 1'h1;
  assign T166 = io_inChannels_1_flit_x[1'h0:1'h0];
  assign T167 = T169 | T168;
  assign T168 = ~ io_inChannels_1_flitValid;
  assign T169 = T170 & T158;
  assign T170 = RouterBuffer_2_io_enq_ready & io_inChannels_1_flitValid;
  assign T172 = T173 | reset;
  assign T173 = T175 | T174;
  assign T174 = T1387 & T158;
  assign T175 = ~ T1387;
  assign T177 = T178 | reset;
  assign T178 = T189 | T179;
  assign T179 = ~ T180;
  assign T180 = T181 == 1'h1;
  assign T181 = T182;
  assign T182 = T187 ? T185 : T183;
  assign T183 = T184[6'h24:6'h24];
  assign T184 = io_inChannels_0_flit_x[6'h36:1'h1];
  assign T185 = T186[4'hd:4'hd];
  assign T186 = io_inChannels_0_flit_x[5'h1f:1'h1];
  assign T187 = T188 == 1'h1;
  assign T188 = io_inChannels_0_flit_x[1'h0:1'h0];
  assign T189 = T191 | T190;
  assign T190 = ~ io_inChannels_0_flitValid;
  assign T191 = T192 & T180;
  assign T192 = RouterBuffer_1_io_enq_ready & io_inChannels_0_flitValid;
  assign T194 = T195 | reset;
  assign T195 = T197 | T196;
  assign T196 = T1531 & T180;
  assign T197 = ~ T1531;
  assign T199 = T200 | reset;
  assign T200 = T211 | T201;
  assign T201 = ~ T202;
  assign T202 = T203 == 1'h0;
  assign T203 = T204;
  assign T204 = T209 ? T207 : T205;
  assign T205 = T206[6'h24:6'h24];
  assign T206 = io_inChannels_0_flit_x[6'h36:1'h1];
  assign T207 = T208[4'hd:4'hd];
  assign T208 = io_inChannels_0_flit_x[5'h1f:1'h1];
  assign T209 = T210 == 1'h1;
  assign T210 = io_inChannels_0_flit_x[1'h0:1'h0];
  assign T211 = T213 | T212;
  assign T212 = ~ io_inChannels_0_flitValid;
  assign T213 = T214 & T202;
  assign T214 = RouterBuffer_io_enq_ready & io_inChannels_0_flitValid;
  assign T216 = T217 | reset;
  assign T217 = T219 | T218;
  assign T218 = T1675 & T202;
  assign T219 = ~ T1675;
  assign T220 = T1722 & T221;
  assign T221 = T222 == 1'h1;
  assign T222 = T223;
  assign T223 = T228 ? T226 : T224;
  assign T224 = T225[6'h24:6'h24];
  assign T225 = switch_io_outPorts_4_x[6'h36:1'h1];
  assign T226 = T227[4'hd:4'hd];
  assign T227 = switch_io_outPorts_4_x[5'h1f:1'h1];
  assign T228 = T229 == 1'h1;
  assign T229 = switch_io_outPorts_4_x[1'h0:1'h0];
  assign T230 = T1722 & T231;
  assign T231 = T222 == 1'h0;
  assign T232 = T1905 & T233;
  assign T233 = T234 == 1'h1;
  assign T234 = T235;
  assign T235 = T240 ? T238 : T236;
  assign T236 = T237[6'h24:6'h24];
  assign T237 = switch_io_outPorts_3_x[6'h36:1'h1];
  assign T238 = T239[4'hd:4'hd];
  assign T239 = switch_io_outPorts_3_x[5'h1f:1'h1];
  assign T240 = T241 == 1'h1;
  assign T241 = switch_io_outPorts_3_x[1'h0:1'h0];
  assign T242 = T1905 & T243;
  assign T243 = T234 == 1'h0;
  assign T244 = T1968 & T245;
  assign T245 = T246 == 1'h1;
  assign T246 = T247;
  assign T247 = T252 ? T250 : T248;
  assign T248 = T249[6'h24:6'h24];
  assign T249 = switch_io_outPorts_2_x[6'h36:1'h1];
  assign T250 = T251[4'hd:4'hd];
  assign T251 = switch_io_outPorts_2_x[5'h1f:1'h1];
  assign T252 = T253 == 1'h1;
  assign T253 = switch_io_outPorts_2_x[1'h0:1'h0];
  assign T254 = T1968 & T255;
  assign T255 = T246 == 1'h0;
  assign T256 = T2031 & T257;
  assign T257 = T258 == 1'h1;
  assign T258 = T259;
  assign T259 = T264 ? T262 : T260;
  assign T260 = T261[6'h24:6'h24];
  assign T261 = switch_io_outPorts_1_x[6'h36:1'h1];
  assign T262 = T263[4'hd:4'hd];
  assign T263 = switch_io_outPorts_1_x[5'h1f:1'h1];
  assign T264 = T265 == 1'h1;
  assign T265 = switch_io_outPorts_1_x[1'h0:1'h0];
  assign T266 = T2031 & T267;
  assign T267 = T258 == 1'h0;
  assign T268 = T2094 & T269;
  assign T269 = T270 == 1'h1;
  assign T270 = T271;
  assign T271 = T276 ? T274 : T272;
  assign T272 = T273[6'h24:6'h24];
  assign T273 = switch_io_outPorts_0_x[6'h36:1'h1];
  assign T274 = T275[4'hd:4'hd];
  assign T275 = switch_io_outPorts_0_x[5'h1f:1'h1];
  assign T276 = T277 == 1'h1;
  assign T277 = switch_io_outPorts_0_x[1'h0:1'h0];
  assign T278 = T2094 & T279;
  assign T279 = T270 == 1'h0;
  assign T280 = T281;
  assign T281 = io_inChannels_4_flit_x;
  assign T3112 = R282[1'h0:1'h0];
  assign T3113 = reset ? 55'h0 : T283;
  assign T283 = T284 ? T3114 : R282;
  assign T3114 = {51'h0, vcAllocator_io_chosens_9};
  assign T284 = T285 & vcAllocator_io_resources_9_valid;
  assign T285 = VCRouterStateManagement_9_io_currentState == 3'h2;
  assign T286 = T287;
  assign T287 = RouterBuffer_9_io_deq_bits_x;
  assign T288 = T300 | T289;
  assign T289 = T290 == 2'h1;
  assign T290 = T299 ? VCRouterOutputStateManagement_4_io_currentState : T291;
  assign T291 = T298 ? T296 : T292;
  assign T292 = T293 ? VCRouterOutputStateManagement_1_io_currentState : VCRouterOutputStateManagement_io_currentState;
  assign T293 = T294[1'h0:1'h0];
  assign T294 = R295;
  assign T3115 = reset ? 3'h0 : CMeshDOR_9_io_result;
  assign T296 = T297 ? VCRouterOutputStateManagement_3_io_currentState : VCRouterOutputStateManagement_2_io_currentState;
  assign T297 = T294[1'h0:1'h0];
  assign T298 = T294[1'h1:1'h1];
  assign T299 = T294[2'h2:2'h2];
  assign T300 = T290 == 2'h2;
  assign T301 = T319 ? T311 : T302;
  assign T302 = T310 ? creditConsReady_4_0 : T303;
  assign T303 = T309 ? T307 : T304;
  assign T304 = T305 ? creditConsReady_1_0 : creditConsReady_0_0;
  assign creditConsReady_0_0 = CreditCon_io_outCredit;
  assign creditConsReady_1_0 = CreditCon_2_io_outCredit;
  assign T305 = T306[1'h0:1'h0];
  assign T306 = R295;
  assign T307 = T308 ? creditConsReady_3_0 : creditConsReady_2_0;
  assign creditConsReady_2_0 = CreditCon_4_io_outCredit;
  assign creditConsReady_3_0 = CreditCon_6_io_outCredit;
  assign T308 = T306[1'h0:1'h0];
  assign T309 = T306[1'h1:1'h1];
  assign creditConsReady_4_0 = CreditCon_8_io_outCredit;
  assign T310 = T306[2'h2:2'h2];
  assign T311 = T318 ? creditConsReady_4_1 : T312;
  assign T312 = T317 ? T315 : T313;
  assign T313 = T314 ? creditConsReady_1_1 : creditConsReady_0_1;
  assign creditConsReady_0_1 = CreditCon_1_io_outCredit;
  assign creditConsReady_1_1 = CreditCon_3_io_outCredit;
  assign T314 = T306[1'h0:1'h0];
  assign T315 = T316 ? creditConsReady_3_1 : creditConsReady_2_1;
  assign creditConsReady_2_1 = CreditCon_5_io_outCredit;
  assign creditConsReady_3_1 = CreditCon_7_io_outCredit;
  assign T316 = T306[1'h0:1'h0];
  assign T317 = T306[1'h1:1'h1];
  assign creditConsReady_4_1 = CreditCon_9_io_outCredit;
  assign T318 = T306[2'h2:2'h2];
  assign T319 = T3116;
  assign T3116 = R282[1'h0:1'h0];
  assign T320 = T331 & T321;
  assign T321 = T322 == 4'h9;
  assign T322 = T330 ? swAllocator_io_chosens_4 : T323;
  assign T323 = T329 ? T327 : T324;
  assign T324 = T325 ? swAllocator_io_chosens_1 : swAllocator_io_chosens_0;
  assign T325 = T326[1'h0:1'h0];
  assign T326 = R295;
  assign T327 = T328 ? swAllocator_io_chosens_3 : swAllocator_io_chosens_2;
  assign T328 = T326[1'h0:1'h0];
  assign T329 = T326[1'h1:1'h1];
  assign T330 = T326[2'h2:2'h2];
  assign T331 = T339 ? swAllocator_io_requests_4_9_grant : T332;
  assign T332 = T338 ? T336 : T333;
  assign T333 = T334 ? swAllocator_io_requests_1_9_grant : swAllocator_io_requests_0_9_grant;
  assign T334 = T335[1'h0:1'h0];
  assign T335 = R295;
  assign T336 = T337 ? swAllocator_io_requests_3_9_grant : swAllocator_io_requests_2_9_grant;
  assign T337 = T335[1'h0:1'h0];
  assign T338 = T335[1'h1:1'h1];
  assign T339 = T335[2'h2:2'h2];
  assign T340 = RouterBuffer_9_io_deq_valid & T341;
  assign T341 = T342;
  assign T342 = T347 ? T345 : T343;
  assign T343 = T344[6'h25:6'h25];
  assign T344 = RouterBuffer_9_io_deq_bits_x[6'h36:1'h1];
  assign T345 = T346[4'he:4'he];
  assign T346 = RouterBuffer_9_io_deq_bits_x[5'h1f:1'h1];
  assign T347 = T348 == 1'h1;
  assign T348 = RouterBuffer_9_io_deq_bits_x[1'h0:1'h0];
  assign T3117 = reset ? 1'h0 : RouterBuffer_9_io_deq_valid;
  assign T350 = T351[2'h2:1'h0];
  assign T351 = T352[5'h1f:1'h1];
  assign T352 = RouterRegFile_9_io_readData;
  assign T353 = T351[3'h4:2'h3];
  assign T354 = T351[3'h6:3'h5];
  assign T355 = T351[4'h8:3'h7];
  assign T356 = T351[4'hc:4'h9];
  assign T357 = T351[4'hd:4'hd];
  assign T358 = T351[4'he:4'he];
  assign T359 = T351[5'h1e:4'hf];
  assign T360 = T374 ? T371 : T361;
  assign T361 = T367 ? 1'h0 : T362;
  assign T362 = T363 & T301;
  assign T363 = T365 & T364;
  assign T364 = VCRouterStateManagement_9_io_currentState == 3'h4;
  assign T365 = T320 | T366;
  assign T366 = VCRouterStateManagement_9_io_currentState == 3'h4;
  assign T367 = T369 & T368;
  assign T368 = ~ RouterRegFile_9_io_readValid;
  assign T369 = T370 == 1'h1;
  assign T370 = RouterBuffer_9_io_deq_bits_x[1'h0:1'h0];
  assign T371 = T372 & T301;
  assign T372 = T365 & T373;
  assign T373 = 3'h3 <= VCRouterStateManagement_9_io_currentState;
  assign T374 = T378 & T375;
  assign T375 = T376 & RouterRegFile_9_io_readValid;
  assign T376 = T377 == 1'h1;
  assign T377 = RouterBuffer_9_io_deq_bits_x[1'h0:1'h0];
  assign T378 = T367 ^ 1'h1;
  assign T379 = io_inChannels_4_flitValid & T4;
  assign T380 = T381 & RouterRegFile_9_io_readValid;
  assign T381 = RouterRegFile_9_io_rvPipelineReg_0 ^ 1'h1;
  assign T382 = T384 & T383;
  assign T383 = VCRouterStateManagement_9_io_currentState == 3'h2;
  assign T384 = RouterRegFile_9_io_rvPipelineReg_0 & vcAllocator_io_resources_9_valid;
  assign T385 = T387 & T386;
  assign T386 = VCRouterStateManagement_9_io_currentState == 3'h3;
  assign T387 = RouterRegFile_9_io_rvPipelineReg_1 & T320;
  assign T3118 = {24'h0, T388};
  assign T388 = T389;
  assign T389 = {T393, T390};
  assign T390 = {T392, T391};
  assign T391 = {CMeshDOR_9_io_outHeadFlit_destination_0, CMeshDOR_9_io_outHeadFlit_priorityLevel};
  assign T392 = {CMeshDOR_9_io_outHeadFlit_destination_2, CMeshDOR_9_io_outHeadFlit_destination_1};
  assign T393 = {T395, T394};
  assign T394 = {CMeshDOR_9_io_outHeadFlit_vcPort, CMeshDOR_9_io_outHeadFlit_packetType};
  assign T395 = {CMeshDOR_9_io_outHeadFlit_packetID, CMeshDOR_9_io_outHeadFlit_isTail};
  assign T396 = T398 & T397;
  assign T397 = VCRouterStateManagement_9_io_currentState == 3'h4;
  assign T398 = T399 & T301;
  assign T399 = T365 & flitsAreTail_9;
  assign flitsAreTail_9 = T400;
  assign T400 = T401 & RouterBuffer_9_io_deq_valid;
  assign T401 = T402;
  assign T402 = T407 ? T405 : T403;
  assign T403 = T404[6'h25:6'h25];
  assign T404 = RouterBuffer_9_io_deq_bits_x[6'h36:1'h1];
  assign T405 = T406[4'he:4'he];
  assign T406 = RouterBuffer_9_io_deq_bits_x[5'h1f:1'h1];
  assign T407 = T408 == 1'h1;
  assign T408 = RouterBuffer_9_io_deq_bits_x[1'h0:1'h0];
  assign T409 = T410 ? T379 : 1'h0;
  assign T410 = T411 == 1'h1;
  assign T411 = io_inChannels_4_flit_x[1'h0:1'h0];
  assign T412 = T410 ? T413 : 55'h0;
  assign T413 = io_inChannels_4_flit_x;
  assign T414 = T374 ? T420 : T415;
  assign T415 = T367 ? 1'h0 : T416;
  assign T416 = T417 & RouterBuffer_9_io_deq_valid;
  assign T417 = T418 & T301;
  assign T418 = T365 & T419;
  assign T419 = VCRouterStateManagement_9_io_currentState == 3'h4;
  assign T420 = T421 & RouterBuffer_9_io_deq_valid;
  assign T421 = T422 & T301;
  assign T422 = T365 & T423;
  assign T423 = 3'h3 <= VCRouterStateManagement_9_io_currentState;
  assign T424 = T425;
  assign T425 = io_inChannels_4_flit_x;
  assign T3119 = R426[1'h0:1'h0];
  assign T3120 = reset ? 55'h0 : T427;
  assign T427 = T428 ? T3121 : R426;
  assign T3121 = {51'h0, vcAllocator_io_chosens_8};
  assign T428 = T429 & vcAllocator_io_resources_8_valid;
  assign T429 = VCRouterStateManagement_8_io_currentState == 3'h2;
  assign T430 = T431;
  assign T431 = RouterBuffer_8_io_deq_bits_x;
  assign T432 = T444 | T433;
  assign T433 = T434 == 2'h1;
  assign T434 = T443 ? VCRouterOutputStateManagement_4_io_currentState : T435;
  assign T435 = T442 ? T440 : T436;
  assign T436 = T437 ? VCRouterOutputStateManagement_1_io_currentState : VCRouterOutputStateManagement_io_currentState;
  assign T437 = T438[1'h0:1'h0];
  assign T438 = R439;
  assign T3122 = reset ? 3'h0 : CMeshDOR_8_io_result;
  assign T440 = T441 ? VCRouterOutputStateManagement_3_io_currentState : VCRouterOutputStateManagement_2_io_currentState;
  assign T441 = T438[1'h0:1'h0];
  assign T442 = T438[1'h1:1'h1];
  assign T443 = T438[2'h2:2'h2];
  assign T444 = T434 == 2'h2;
  assign T445 = T463 ? T455 : T446;
  assign T446 = T454 ? creditConsReady_4_0 : T447;
  assign T447 = T453 ? T451 : T448;
  assign T448 = T449 ? creditConsReady_1_0 : creditConsReady_0_0;
  assign T449 = T450[1'h0:1'h0];
  assign T450 = R439;
  assign T451 = T452 ? creditConsReady_3_0 : creditConsReady_2_0;
  assign T452 = T450[1'h0:1'h0];
  assign T453 = T450[1'h1:1'h1];
  assign T454 = T450[2'h2:2'h2];
  assign T455 = T462 ? creditConsReady_4_1 : T456;
  assign T456 = T461 ? T459 : T457;
  assign T457 = T458 ? creditConsReady_1_1 : creditConsReady_0_1;
  assign T458 = T450[1'h0:1'h0];
  assign T459 = T460 ? creditConsReady_3_1 : creditConsReady_2_1;
  assign T460 = T450[1'h0:1'h0];
  assign T461 = T450[1'h1:1'h1];
  assign T462 = T450[2'h2:2'h2];
  assign T463 = T3123;
  assign T3123 = R426[1'h0:1'h0];
  assign T464 = T475 & T465;
  assign T465 = T466 == 4'h8;
  assign T466 = T474 ? swAllocator_io_chosens_4 : T467;
  assign T467 = T473 ? T471 : T468;
  assign T468 = T469 ? swAllocator_io_chosens_1 : swAllocator_io_chosens_0;
  assign T469 = T470[1'h0:1'h0];
  assign T470 = R439;
  assign T471 = T472 ? swAllocator_io_chosens_3 : swAllocator_io_chosens_2;
  assign T472 = T470[1'h0:1'h0];
  assign T473 = T470[1'h1:1'h1];
  assign T474 = T470[2'h2:2'h2];
  assign T475 = T483 ? swAllocator_io_requests_4_8_grant : T476;
  assign T476 = T482 ? T480 : T477;
  assign T477 = T478 ? swAllocator_io_requests_1_8_grant : swAllocator_io_requests_0_8_grant;
  assign T478 = T479[1'h0:1'h0];
  assign T479 = R439;
  assign T480 = T481 ? swAllocator_io_requests_3_8_grant : swAllocator_io_requests_2_8_grant;
  assign T481 = T479[1'h0:1'h0];
  assign T482 = T479[1'h1:1'h1];
  assign T483 = T479[2'h2:2'h2];
  assign T484 = RouterBuffer_8_io_deq_valid & T485;
  assign T485 = T486;
  assign T486 = T491 ? T489 : T487;
  assign T487 = T488[6'h25:6'h25];
  assign T488 = RouterBuffer_8_io_deq_bits_x[6'h36:1'h1];
  assign T489 = T490[4'he:4'he];
  assign T490 = RouterBuffer_8_io_deq_bits_x[5'h1f:1'h1];
  assign T491 = T492 == 1'h1;
  assign T492 = RouterBuffer_8_io_deq_bits_x[1'h0:1'h0];
  assign T3124 = reset ? 1'h0 : RouterBuffer_8_io_deq_valid;
  assign T494 = T495[2'h2:1'h0];
  assign T495 = T496[5'h1f:1'h1];
  assign T496 = RouterRegFile_8_io_readData;
  assign T497 = T495[3'h4:2'h3];
  assign T498 = T495[3'h6:3'h5];
  assign T499 = T495[4'h8:3'h7];
  assign T500 = T495[4'hc:4'h9];
  assign T501 = T495[4'hd:4'hd];
  assign T502 = T495[4'he:4'he];
  assign T503 = T495[5'h1e:4'hf];
  assign T504 = T518 ? T515 : T505;
  assign T505 = T511 ? 1'h0 : T506;
  assign T506 = T507 & T445;
  assign T507 = T509 & T508;
  assign T508 = VCRouterStateManagement_8_io_currentState == 3'h4;
  assign T509 = T464 | T510;
  assign T510 = VCRouterStateManagement_8_io_currentState == 3'h4;
  assign T511 = T513 & T512;
  assign T512 = ~ RouterRegFile_8_io_readValid;
  assign T513 = T514 == 1'h1;
  assign T514 = RouterBuffer_8_io_deq_bits_x[1'h0:1'h0];
  assign T515 = T516 & T445;
  assign T516 = T509 & T517;
  assign T517 = 3'h3 <= VCRouterStateManagement_8_io_currentState;
  assign T518 = T522 & T519;
  assign T519 = T520 & RouterRegFile_8_io_readValid;
  assign T520 = T521 == 1'h1;
  assign T521 = RouterBuffer_8_io_deq_bits_x[1'h0:1'h0];
  assign T522 = T511 ^ 1'h1;
  assign T523 = io_inChannels_4_flitValid & T26;
  assign T524 = T525 & RouterRegFile_8_io_readValid;
  assign T525 = RouterRegFile_8_io_rvPipelineReg_0 ^ 1'h1;
  assign T526 = T528 & T527;
  assign T527 = VCRouterStateManagement_8_io_currentState == 3'h2;
  assign T528 = RouterRegFile_8_io_rvPipelineReg_0 & vcAllocator_io_resources_8_valid;
  assign T529 = T531 & T530;
  assign T530 = VCRouterStateManagement_8_io_currentState == 3'h3;
  assign T531 = RouterRegFile_8_io_rvPipelineReg_1 & T464;
  assign T3125 = {24'h0, T532};
  assign T532 = T533;
  assign T533 = {T537, T534};
  assign T534 = {T536, T535};
  assign T535 = {CMeshDOR_8_io_outHeadFlit_destination_0, CMeshDOR_8_io_outHeadFlit_priorityLevel};
  assign T536 = {CMeshDOR_8_io_outHeadFlit_destination_2, CMeshDOR_8_io_outHeadFlit_destination_1};
  assign T537 = {T539, T538};
  assign T538 = {CMeshDOR_8_io_outHeadFlit_vcPort, CMeshDOR_8_io_outHeadFlit_packetType};
  assign T539 = {CMeshDOR_8_io_outHeadFlit_packetID, CMeshDOR_8_io_outHeadFlit_isTail};
  assign T540 = T542 & T541;
  assign T541 = VCRouterStateManagement_8_io_currentState == 3'h4;
  assign T542 = T543 & T445;
  assign T543 = T509 & flitsAreTail_8;
  assign flitsAreTail_8 = T544;
  assign T544 = T545 & RouterBuffer_8_io_deq_valid;
  assign T545 = T546;
  assign T546 = T551 ? T549 : T547;
  assign T547 = T548[6'h25:6'h25];
  assign T548 = RouterBuffer_8_io_deq_bits_x[6'h36:1'h1];
  assign T549 = T550[4'he:4'he];
  assign T550 = RouterBuffer_8_io_deq_bits_x[5'h1f:1'h1];
  assign T551 = T552 == 1'h1;
  assign T552 = RouterBuffer_8_io_deq_bits_x[1'h0:1'h0];
  assign T553 = T554 ? T523 : 1'h0;
  assign T554 = T555 == 1'h1;
  assign T555 = io_inChannels_4_flit_x[1'h0:1'h0];
  assign T556 = T554 ? T557 : 55'h0;
  assign T557 = io_inChannels_4_flit_x;
  assign T558 = T518 ? T564 : T559;
  assign T559 = T511 ? 1'h0 : T560;
  assign T560 = T561 & RouterBuffer_8_io_deq_valid;
  assign T561 = T562 & T445;
  assign T562 = T509 & T563;
  assign T563 = VCRouterStateManagement_8_io_currentState == 3'h4;
  assign T564 = T565 & RouterBuffer_8_io_deq_valid;
  assign T565 = T566 & T445;
  assign T566 = T509 & T567;
  assign T567 = 3'h3 <= VCRouterStateManagement_8_io_currentState;
  assign T568 = T569;
  assign T569 = io_inChannels_3_flit_x;
  assign T3126 = R570[1'h0:1'h0];
  assign T3127 = reset ? 55'h0 : T571;
  assign T571 = T572 ? T3128 : R570;
  assign T3128 = {51'h0, vcAllocator_io_chosens_7};
  assign T572 = T573 & vcAllocator_io_resources_7_valid;
  assign T573 = VCRouterStateManagement_7_io_currentState == 3'h2;
  assign T574 = T575;
  assign T575 = RouterBuffer_7_io_deq_bits_x;
  assign T576 = T588 | T577;
  assign T577 = T578 == 2'h1;
  assign T578 = T587 ? VCRouterOutputStateManagement_4_io_currentState : T579;
  assign T579 = T586 ? T584 : T580;
  assign T580 = T581 ? VCRouterOutputStateManagement_1_io_currentState : VCRouterOutputStateManagement_io_currentState;
  assign T581 = T582[1'h0:1'h0];
  assign T582 = R583;
  assign T3129 = reset ? 3'h0 : CMeshDOR_7_io_result;
  assign T584 = T585 ? VCRouterOutputStateManagement_3_io_currentState : VCRouterOutputStateManagement_2_io_currentState;
  assign T585 = T582[1'h0:1'h0];
  assign T586 = T582[1'h1:1'h1];
  assign T587 = T582[2'h2:2'h2];
  assign T588 = T578 == 2'h2;
  assign T589 = T607 ? T599 : T590;
  assign T590 = T598 ? creditConsReady_4_0 : T591;
  assign T591 = T597 ? T595 : T592;
  assign T592 = T593 ? creditConsReady_1_0 : creditConsReady_0_0;
  assign T593 = T594[1'h0:1'h0];
  assign T594 = R583;
  assign T595 = T596 ? creditConsReady_3_0 : creditConsReady_2_0;
  assign T596 = T594[1'h0:1'h0];
  assign T597 = T594[1'h1:1'h1];
  assign T598 = T594[2'h2:2'h2];
  assign T599 = T606 ? creditConsReady_4_1 : T600;
  assign T600 = T605 ? T603 : T601;
  assign T601 = T602 ? creditConsReady_1_1 : creditConsReady_0_1;
  assign T602 = T594[1'h0:1'h0];
  assign T603 = T604 ? creditConsReady_3_1 : creditConsReady_2_1;
  assign T604 = T594[1'h0:1'h0];
  assign T605 = T594[1'h1:1'h1];
  assign T606 = T594[2'h2:2'h2];
  assign T607 = T3130;
  assign T3130 = R570[1'h0:1'h0];
  assign T608 = T619 & T609;
  assign T609 = T610 == 4'h7;
  assign T610 = T618 ? swAllocator_io_chosens_4 : T611;
  assign T611 = T617 ? T615 : T612;
  assign T612 = T613 ? swAllocator_io_chosens_1 : swAllocator_io_chosens_0;
  assign T613 = T614[1'h0:1'h0];
  assign T614 = R583;
  assign T615 = T616 ? swAllocator_io_chosens_3 : swAllocator_io_chosens_2;
  assign T616 = T614[1'h0:1'h0];
  assign T617 = T614[1'h1:1'h1];
  assign T618 = T614[2'h2:2'h2];
  assign T619 = T627 ? swAllocator_io_requests_4_7_grant : T620;
  assign T620 = T626 ? T624 : T621;
  assign T621 = T622 ? swAllocator_io_requests_1_7_grant : swAllocator_io_requests_0_7_grant;
  assign T622 = T623[1'h0:1'h0];
  assign T623 = R583;
  assign T624 = T625 ? swAllocator_io_requests_3_7_grant : swAllocator_io_requests_2_7_grant;
  assign T625 = T623[1'h0:1'h0];
  assign T626 = T623[1'h1:1'h1];
  assign T627 = T623[2'h2:2'h2];
  assign T628 = RouterBuffer_7_io_deq_valid & T629;
  assign T629 = T630;
  assign T630 = T635 ? T633 : T631;
  assign T631 = T632[6'h25:6'h25];
  assign T632 = RouterBuffer_7_io_deq_bits_x[6'h36:1'h1];
  assign T633 = T634[4'he:4'he];
  assign T634 = RouterBuffer_7_io_deq_bits_x[5'h1f:1'h1];
  assign T635 = T636 == 1'h1;
  assign T636 = RouterBuffer_7_io_deq_bits_x[1'h0:1'h0];
  assign T3131 = reset ? 1'h0 : RouterBuffer_7_io_deq_valid;
  assign T638 = T639[2'h2:1'h0];
  assign T639 = T640[5'h1f:1'h1];
  assign T640 = RouterRegFile_7_io_readData;
  assign T641 = T639[3'h4:2'h3];
  assign T642 = T639[3'h6:3'h5];
  assign T643 = T639[4'h8:3'h7];
  assign T644 = T639[4'hc:4'h9];
  assign T645 = T639[4'hd:4'hd];
  assign T646 = T639[4'he:4'he];
  assign T647 = T639[5'h1e:4'hf];
  assign T648 = T662 ? T659 : T649;
  assign T649 = T655 ? 1'h0 : T650;
  assign T650 = T651 & T589;
  assign T651 = T653 & T652;
  assign T652 = VCRouterStateManagement_7_io_currentState == 3'h4;
  assign T653 = T608 | T654;
  assign T654 = VCRouterStateManagement_7_io_currentState == 3'h4;
  assign T655 = T657 & T656;
  assign T656 = ~ RouterRegFile_7_io_readValid;
  assign T657 = T658 == 1'h1;
  assign T658 = RouterBuffer_7_io_deq_bits_x[1'h0:1'h0];
  assign T659 = T660 & T589;
  assign T660 = T653 & T661;
  assign T661 = 3'h3 <= VCRouterStateManagement_7_io_currentState;
  assign T662 = T666 & T663;
  assign T663 = T664 & RouterRegFile_7_io_readValid;
  assign T664 = T665 == 1'h1;
  assign T665 = RouterBuffer_7_io_deq_bits_x[1'h0:1'h0];
  assign T666 = T655 ^ 1'h1;
  assign T667 = io_inChannels_3_flitValid & T48;
  assign T668 = T669 & RouterRegFile_7_io_readValid;
  assign T669 = RouterRegFile_7_io_rvPipelineReg_0 ^ 1'h1;
  assign T670 = T672 & T671;
  assign T671 = VCRouterStateManagement_7_io_currentState == 3'h2;
  assign T672 = RouterRegFile_7_io_rvPipelineReg_0 & vcAllocator_io_resources_7_valid;
  assign T673 = T675 & T674;
  assign T674 = VCRouterStateManagement_7_io_currentState == 3'h3;
  assign T675 = RouterRegFile_7_io_rvPipelineReg_1 & T608;
  assign T3132 = {24'h0, T676};
  assign T676 = T677;
  assign T677 = {T681, T678};
  assign T678 = {T680, T679};
  assign T679 = {CMeshDOR_7_io_outHeadFlit_destination_0, CMeshDOR_7_io_outHeadFlit_priorityLevel};
  assign T680 = {CMeshDOR_7_io_outHeadFlit_destination_2, CMeshDOR_7_io_outHeadFlit_destination_1};
  assign T681 = {T683, T682};
  assign T682 = {CMeshDOR_7_io_outHeadFlit_vcPort, CMeshDOR_7_io_outHeadFlit_packetType};
  assign T683 = {CMeshDOR_7_io_outHeadFlit_packetID, CMeshDOR_7_io_outHeadFlit_isTail};
  assign T684 = T686 & T685;
  assign T685 = VCRouterStateManagement_7_io_currentState == 3'h4;
  assign T686 = T687 & T589;
  assign T687 = T653 & flitsAreTail_7;
  assign flitsAreTail_7 = T688;
  assign T688 = T689 & RouterBuffer_7_io_deq_valid;
  assign T689 = T690;
  assign T690 = T695 ? T693 : T691;
  assign T691 = T692[6'h25:6'h25];
  assign T692 = RouterBuffer_7_io_deq_bits_x[6'h36:1'h1];
  assign T693 = T694[4'he:4'he];
  assign T694 = RouterBuffer_7_io_deq_bits_x[5'h1f:1'h1];
  assign T695 = T696 == 1'h1;
  assign T696 = RouterBuffer_7_io_deq_bits_x[1'h0:1'h0];
  assign T697 = T698 ? T667 : 1'h0;
  assign T698 = T699 == 1'h1;
  assign T699 = io_inChannels_3_flit_x[1'h0:1'h0];
  assign T700 = T698 ? T701 : 55'h0;
  assign T701 = io_inChannels_3_flit_x;
  assign T702 = T662 ? T708 : T703;
  assign T703 = T655 ? 1'h0 : T704;
  assign T704 = T705 & RouterBuffer_7_io_deq_valid;
  assign T705 = T706 & T589;
  assign T706 = T653 & T707;
  assign T707 = VCRouterStateManagement_7_io_currentState == 3'h4;
  assign T708 = T709 & RouterBuffer_7_io_deq_valid;
  assign T709 = T710 & T589;
  assign T710 = T653 & T711;
  assign T711 = 3'h3 <= VCRouterStateManagement_7_io_currentState;
  assign T712 = T713;
  assign T713 = io_inChannels_3_flit_x;
  assign T3133 = R714[1'h0:1'h0];
  assign T3134 = reset ? 55'h0 : T715;
  assign T715 = T716 ? T3135 : R714;
  assign T3135 = {51'h0, vcAllocator_io_chosens_6};
  assign T716 = T717 & vcAllocator_io_resources_6_valid;
  assign T717 = VCRouterStateManagement_6_io_currentState == 3'h2;
  assign T718 = T719;
  assign T719 = RouterBuffer_6_io_deq_bits_x;
  assign T720 = T732 | T721;
  assign T721 = T722 == 2'h1;
  assign T722 = T731 ? VCRouterOutputStateManagement_4_io_currentState : T723;
  assign T723 = T730 ? T728 : T724;
  assign T724 = T725 ? VCRouterOutputStateManagement_1_io_currentState : VCRouterOutputStateManagement_io_currentState;
  assign T725 = T726[1'h0:1'h0];
  assign T726 = R727;
  assign T3136 = reset ? 3'h0 : CMeshDOR_6_io_result;
  assign T728 = T729 ? VCRouterOutputStateManagement_3_io_currentState : VCRouterOutputStateManagement_2_io_currentState;
  assign T729 = T726[1'h0:1'h0];
  assign T730 = T726[1'h1:1'h1];
  assign T731 = T726[2'h2:2'h2];
  assign T732 = T722 == 2'h2;
  assign T733 = T751 ? T743 : T734;
  assign T734 = T742 ? creditConsReady_4_0 : T735;
  assign T735 = T741 ? T739 : T736;
  assign T736 = T737 ? creditConsReady_1_0 : creditConsReady_0_0;
  assign T737 = T738[1'h0:1'h0];
  assign T738 = R727;
  assign T739 = T740 ? creditConsReady_3_0 : creditConsReady_2_0;
  assign T740 = T738[1'h0:1'h0];
  assign T741 = T738[1'h1:1'h1];
  assign T742 = T738[2'h2:2'h2];
  assign T743 = T750 ? creditConsReady_4_1 : T744;
  assign T744 = T749 ? T747 : T745;
  assign T745 = T746 ? creditConsReady_1_1 : creditConsReady_0_1;
  assign T746 = T738[1'h0:1'h0];
  assign T747 = T748 ? creditConsReady_3_1 : creditConsReady_2_1;
  assign T748 = T738[1'h0:1'h0];
  assign T749 = T738[1'h1:1'h1];
  assign T750 = T738[2'h2:2'h2];
  assign T751 = T3137;
  assign T3137 = R714[1'h0:1'h0];
  assign T752 = T763 & T753;
  assign T753 = T754 == 4'h6;
  assign T754 = T762 ? swAllocator_io_chosens_4 : T755;
  assign T755 = T761 ? T759 : T756;
  assign T756 = T757 ? swAllocator_io_chosens_1 : swAllocator_io_chosens_0;
  assign T757 = T758[1'h0:1'h0];
  assign T758 = R727;
  assign T759 = T760 ? swAllocator_io_chosens_3 : swAllocator_io_chosens_2;
  assign T760 = T758[1'h0:1'h0];
  assign T761 = T758[1'h1:1'h1];
  assign T762 = T758[2'h2:2'h2];
  assign T763 = T771 ? swAllocator_io_requests_4_6_grant : T764;
  assign T764 = T770 ? T768 : T765;
  assign T765 = T766 ? swAllocator_io_requests_1_6_grant : swAllocator_io_requests_0_6_grant;
  assign T766 = T767[1'h0:1'h0];
  assign T767 = R727;
  assign T768 = T769 ? swAllocator_io_requests_3_6_grant : swAllocator_io_requests_2_6_grant;
  assign T769 = T767[1'h0:1'h0];
  assign T770 = T767[1'h1:1'h1];
  assign T771 = T767[2'h2:2'h2];
  assign T772 = RouterBuffer_6_io_deq_valid & T773;
  assign T773 = T774;
  assign T774 = T779 ? T777 : T775;
  assign T775 = T776[6'h25:6'h25];
  assign T776 = RouterBuffer_6_io_deq_bits_x[6'h36:1'h1];
  assign T777 = T778[4'he:4'he];
  assign T778 = RouterBuffer_6_io_deq_bits_x[5'h1f:1'h1];
  assign T779 = T780 == 1'h1;
  assign T780 = RouterBuffer_6_io_deq_bits_x[1'h0:1'h0];
  assign T3138 = reset ? 1'h0 : RouterBuffer_6_io_deq_valid;
  assign T782 = T783[2'h2:1'h0];
  assign T783 = T784[5'h1f:1'h1];
  assign T784 = RouterRegFile_6_io_readData;
  assign T785 = T783[3'h4:2'h3];
  assign T786 = T783[3'h6:3'h5];
  assign T787 = T783[4'h8:3'h7];
  assign T788 = T783[4'hc:4'h9];
  assign T789 = T783[4'hd:4'hd];
  assign T790 = T783[4'he:4'he];
  assign T791 = T783[5'h1e:4'hf];
  assign T792 = T806 ? T803 : T793;
  assign T793 = T799 ? 1'h0 : T794;
  assign T794 = T795 & T733;
  assign T795 = T797 & T796;
  assign T796 = VCRouterStateManagement_6_io_currentState == 3'h4;
  assign T797 = T752 | T798;
  assign T798 = VCRouterStateManagement_6_io_currentState == 3'h4;
  assign T799 = T801 & T800;
  assign T800 = ~ RouterRegFile_6_io_readValid;
  assign T801 = T802 == 1'h1;
  assign T802 = RouterBuffer_6_io_deq_bits_x[1'h0:1'h0];
  assign T803 = T804 & T733;
  assign T804 = T797 & T805;
  assign T805 = 3'h3 <= VCRouterStateManagement_6_io_currentState;
  assign T806 = T810 & T807;
  assign T807 = T808 & RouterRegFile_6_io_readValid;
  assign T808 = T809 == 1'h1;
  assign T809 = RouterBuffer_6_io_deq_bits_x[1'h0:1'h0];
  assign T810 = T799 ^ 1'h1;
  assign T811 = io_inChannels_3_flitValid & T70;
  assign T812 = T813 & RouterRegFile_6_io_readValid;
  assign T813 = RouterRegFile_6_io_rvPipelineReg_0 ^ 1'h1;
  assign T814 = T816 & T815;
  assign T815 = VCRouterStateManagement_6_io_currentState == 3'h2;
  assign T816 = RouterRegFile_6_io_rvPipelineReg_0 & vcAllocator_io_resources_6_valid;
  assign T817 = T819 & T818;
  assign T818 = VCRouterStateManagement_6_io_currentState == 3'h3;
  assign T819 = RouterRegFile_6_io_rvPipelineReg_1 & T752;
  assign T3139 = {24'h0, T820};
  assign T820 = T821;
  assign T821 = {T825, T822};
  assign T822 = {T824, T823};
  assign T823 = {CMeshDOR_6_io_outHeadFlit_destination_0, CMeshDOR_6_io_outHeadFlit_priorityLevel};
  assign T824 = {CMeshDOR_6_io_outHeadFlit_destination_2, CMeshDOR_6_io_outHeadFlit_destination_1};
  assign T825 = {T827, T826};
  assign T826 = {CMeshDOR_6_io_outHeadFlit_vcPort, CMeshDOR_6_io_outHeadFlit_packetType};
  assign T827 = {CMeshDOR_6_io_outHeadFlit_packetID, CMeshDOR_6_io_outHeadFlit_isTail};
  assign T828 = T830 & T829;
  assign T829 = VCRouterStateManagement_6_io_currentState == 3'h4;
  assign T830 = T831 & T733;
  assign T831 = T797 & flitsAreTail_6;
  assign flitsAreTail_6 = T832;
  assign T832 = T833 & RouterBuffer_6_io_deq_valid;
  assign T833 = T834;
  assign T834 = T839 ? T837 : T835;
  assign T835 = T836[6'h25:6'h25];
  assign T836 = RouterBuffer_6_io_deq_bits_x[6'h36:1'h1];
  assign T837 = T838[4'he:4'he];
  assign T838 = RouterBuffer_6_io_deq_bits_x[5'h1f:1'h1];
  assign T839 = T840 == 1'h1;
  assign T840 = RouterBuffer_6_io_deq_bits_x[1'h0:1'h0];
  assign T841 = T842 ? T811 : 1'h0;
  assign T842 = T843 == 1'h1;
  assign T843 = io_inChannels_3_flit_x[1'h0:1'h0];
  assign T844 = T842 ? T845 : 55'h0;
  assign T845 = io_inChannels_3_flit_x;
  assign T846 = T806 ? T852 : T847;
  assign T847 = T799 ? 1'h0 : T848;
  assign T848 = T849 & RouterBuffer_6_io_deq_valid;
  assign T849 = T850 & T733;
  assign T850 = T797 & T851;
  assign T851 = VCRouterStateManagement_6_io_currentState == 3'h4;
  assign T852 = T853 & RouterBuffer_6_io_deq_valid;
  assign T853 = T854 & T733;
  assign T854 = T797 & T855;
  assign T855 = 3'h3 <= VCRouterStateManagement_6_io_currentState;
  assign T856 = T857;
  assign T857 = io_inChannels_2_flit_x;
  assign T3140 = R858[1'h0:1'h0];
  assign T3141 = reset ? 55'h0 : T859;
  assign T859 = T860 ? T3142 : R858;
  assign T3142 = {51'h0, vcAllocator_io_chosens_5};
  assign T860 = T861 & vcAllocator_io_resources_5_valid;
  assign T861 = VCRouterStateManagement_5_io_currentState == 3'h2;
  assign T862 = T863;
  assign T863 = RouterBuffer_5_io_deq_bits_x;
  assign T864 = T876 | T865;
  assign T865 = T866 == 2'h1;
  assign T866 = T875 ? VCRouterOutputStateManagement_4_io_currentState : T867;
  assign T867 = T874 ? T872 : T868;
  assign T868 = T869 ? VCRouterOutputStateManagement_1_io_currentState : VCRouterOutputStateManagement_io_currentState;
  assign T869 = T870[1'h0:1'h0];
  assign T870 = R871;
  assign T3143 = reset ? 3'h0 : CMeshDOR_5_io_result;
  assign T872 = T873 ? VCRouterOutputStateManagement_3_io_currentState : VCRouterOutputStateManagement_2_io_currentState;
  assign T873 = T870[1'h0:1'h0];
  assign T874 = T870[1'h1:1'h1];
  assign T875 = T870[2'h2:2'h2];
  assign T876 = T866 == 2'h2;
  assign T877 = T895 ? T887 : T878;
  assign T878 = T886 ? creditConsReady_4_0 : T879;
  assign T879 = T885 ? T883 : T880;
  assign T880 = T881 ? creditConsReady_1_0 : creditConsReady_0_0;
  assign T881 = T882[1'h0:1'h0];
  assign T882 = R871;
  assign T883 = T884 ? creditConsReady_3_0 : creditConsReady_2_0;
  assign T884 = T882[1'h0:1'h0];
  assign T885 = T882[1'h1:1'h1];
  assign T886 = T882[2'h2:2'h2];
  assign T887 = T894 ? creditConsReady_4_1 : T888;
  assign T888 = T893 ? T891 : T889;
  assign T889 = T890 ? creditConsReady_1_1 : creditConsReady_0_1;
  assign T890 = T882[1'h0:1'h0];
  assign T891 = T892 ? creditConsReady_3_1 : creditConsReady_2_1;
  assign T892 = T882[1'h0:1'h0];
  assign T893 = T882[1'h1:1'h1];
  assign T894 = T882[2'h2:2'h2];
  assign T895 = T3144;
  assign T3144 = R858[1'h0:1'h0];
  assign T896 = T907 & T897;
  assign T897 = T898 == 4'h5;
  assign T898 = T906 ? swAllocator_io_chosens_4 : T899;
  assign T899 = T905 ? T903 : T900;
  assign T900 = T901 ? swAllocator_io_chosens_1 : swAllocator_io_chosens_0;
  assign T901 = T902[1'h0:1'h0];
  assign T902 = R871;
  assign T903 = T904 ? swAllocator_io_chosens_3 : swAllocator_io_chosens_2;
  assign T904 = T902[1'h0:1'h0];
  assign T905 = T902[1'h1:1'h1];
  assign T906 = T902[2'h2:2'h2];
  assign T907 = T915 ? swAllocator_io_requests_4_5_grant : T908;
  assign T908 = T914 ? T912 : T909;
  assign T909 = T910 ? swAllocator_io_requests_1_5_grant : swAllocator_io_requests_0_5_grant;
  assign T910 = T911[1'h0:1'h0];
  assign T911 = R871;
  assign T912 = T913 ? swAllocator_io_requests_3_5_grant : swAllocator_io_requests_2_5_grant;
  assign T913 = T911[1'h0:1'h0];
  assign T914 = T911[1'h1:1'h1];
  assign T915 = T911[2'h2:2'h2];
  assign T916 = RouterBuffer_5_io_deq_valid & T917;
  assign T917 = T918;
  assign T918 = T923 ? T921 : T919;
  assign T919 = T920[6'h25:6'h25];
  assign T920 = RouterBuffer_5_io_deq_bits_x[6'h36:1'h1];
  assign T921 = T922[4'he:4'he];
  assign T922 = RouterBuffer_5_io_deq_bits_x[5'h1f:1'h1];
  assign T923 = T924 == 1'h1;
  assign T924 = RouterBuffer_5_io_deq_bits_x[1'h0:1'h0];
  assign T3145 = reset ? 1'h0 : RouterBuffer_5_io_deq_valid;
  assign T926 = T927[2'h2:1'h0];
  assign T927 = T928[5'h1f:1'h1];
  assign T928 = RouterRegFile_5_io_readData;
  assign T929 = T927[3'h4:2'h3];
  assign T930 = T927[3'h6:3'h5];
  assign T931 = T927[4'h8:3'h7];
  assign T932 = T927[4'hc:4'h9];
  assign T933 = T927[4'hd:4'hd];
  assign T934 = T927[4'he:4'he];
  assign T935 = T927[5'h1e:4'hf];
  assign T936 = T950 ? T947 : T937;
  assign T937 = T943 ? 1'h0 : T938;
  assign T938 = T939 & T877;
  assign T939 = T941 & T940;
  assign T940 = VCRouterStateManagement_5_io_currentState == 3'h4;
  assign T941 = T896 | T942;
  assign T942 = VCRouterStateManagement_5_io_currentState == 3'h4;
  assign T943 = T945 & T944;
  assign T944 = ~ RouterRegFile_5_io_readValid;
  assign T945 = T946 == 1'h1;
  assign T946 = RouterBuffer_5_io_deq_bits_x[1'h0:1'h0];
  assign T947 = T948 & T877;
  assign T948 = T941 & T949;
  assign T949 = 3'h3 <= VCRouterStateManagement_5_io_currentState;
  assign T950 = T954 & T951;
  assign T951 = T952 & RouterRegFile_5_io_readValid;
  assign T952 = T953 == 1'h1;
  assign T953 = RouterBuffer_5_io_deq_bits_x[1'h0:1'h0];
  assign T954 = T943 ^ 1'h1;
  assign T955 = io_inChannels_2_flitValid & T92;
  assign T956 = T957 & RouterRegFile_5_io_readValid;
  assign T957 = RouterRegFile_5_io_rvPipelineReg_0 ^ 1'h1;
  assign T958 = T960 & T959;
  assign T959 = VCRouterStateManagement_5_io_currentState == 3'h2;
  assign T960 = RouterRegFile_5_io_rvPipelineReg_0 & vcAllocator_io_resources_5_valid;
  assign T961 = T963 & T962;
  assign T962 = VCRouterStateManagement_5_io_currentState == 3'h3;
  assign T963 = RouterRegFile_5_io_rvPipelineReg_1 & T896;
  assign T3146 = {24'h0, T964};
  assign T964 = T965;
  assign T965 = {T969, T966};
  assign T966 = {T968, T967};
  assign T967 = {CMeshDOR_5_io_outHeadFlit_destination_0, CMeshDOR_5_io_outHeadFlit_priorityLevel};
  assign T968 = {CMeshDOR_5_io_outHeadFlit_destination_2, CMeshDOR_5_io_outHeadFlit_destination_1};
  assign T969 = {T971, T970};
  assign T970 = {CMeshDOR_5_io_outHeadFlit_vcPort, CMeshDOR_5_io_outHeadFlit_packetType};
  assign T971 = {CMeshDOR_5_io_outHeadFlit_packetID, CMeshDOR_5_io_outHeadFlit_isTail};
  assign T972 = T974 & T973;
  assign T973 = VCRouterStateManagement_5_io_currentState == 3'h4;
  assign T974 = T975 & T877;
  assign T975 = T941 & flitsAreTail_5;
  assign flitsAreTail_5 = T976;
  assign T976 = T977 & RouterBuffer_5_io_deq_valid;
  assign T977 = T978;
  assign T978 = T983 ? T981 : T979;
  assign T979 = T980[6'h25:6'h25];
  assign T980 = RouterBuffer_5_io_deq_bits_x[6'h36:1'h1];
  assign T981 = T982[4'he:4'he];
  assign T982 = RouterBuffer_5_io_deq_bits_x[5'h1f:1'h1];
  assign T983 = T984 == 1'h1;
  assign T984 = RouterBuffer_5_io_deq_bits_x[1'h0:1'h0];
  assign T985 = T986 ? T955 : 1'h0;
  assign T986 = T987 == 1'h1;
  assign T987 = io_inChannels_2_flit_x[1'h0:1'h0];
  assign T988 = T986 ? T989 : 55'h0;
  assign T989 = io_inChannels_2_flit_x;
  assign T990 = T950 ? T996 : T991;
  assign T991 = T943 ? 1'h0 : T992;
  assign T992 = T993 & RouterBuffer_5_io_deq_valid;
  assign T993 = T994 & T877;
  assign T994 = T941 & T995;
  assign T995 = VCRouterStateManagement_5_io_currentState == 3'h4;
  assign T996 = T997 & RouterBuffer_5_io_deq_valid;
  assign T997 = T998 & T877;
  assign T998 = T941 & T999;
  assign T999 = 3'h3 <= VCRouterStateManagement_5_io_currentState;
  assign T1000 = T1001;
  assign T1001 = io_inChannels_2_flit_x;
  assign T3147 = R1002[1'h0:1'h0];
  assign T3148 = reset ? 55'h0 : T1003;
  assign T1003 = T1004 ? T3149 : R1002;
  assign T3149 = {51'h0, vcAllocator_io_chosens_4};
  assign T1004 = T1005 & vcAllocator_io_resources_4_valid;
  assign T1005 = VCRouterStateManagement_4_io_currentState == 3'h2;
  assign T1006 = T1007;
  assign T1007 = RouterBuffer_4_io_deq_bits_x;
  assign T1008 = T1020 | T1009;
  assign T1009 = T1010 == 2'h1;
  assign T1010 = T1019 ? VCRouterOutputStateManagement_4_io_currentState : T1011;
  assign T1011 = T1018 ? T1016 : T1012;
  assign T1012 = T1013 ? VCRouterOutputStateManagement_1_io_currentState : VCRouterOutputStateManagement_io_currentState;
  assign T1013 = T1014[1'h0:1'h0];
  assign T1014 = R1015;
  assign T3150 = reset ? 3'h0 : CMeshDOR_4_io_result;
  assign T1016 = T1017 ? VCRouterOutputStateManagement_3_io_currentState : VCRouterOutputStateManagement_2_io_currentState;
  assign T1017 = T1014[1'h0:1'h0];
  assign T1018 = T1014[1'h1:1'h1];
  assign T1019 = T1014[2'h2:2'h2];
  assign T1020 = T1010 == 2'h2;
  assign T1021 = T1039 ? T1031 : T1022;
  assign T1022 = T1030 ? creditConsReady_4_0 : T1023;
  assign T1023 = T1029 ? T1027 : T1024;
  assign T1024 = T1025 ? creditConsReady_1_0 : creditConsReady_0_0;
  assign T1025 = T1026[1'h0:1'h0];
  assign T1026 = R1015;
  assign T1027 = T1028 ? creditConsReady_3_0 : creditConsReady_2_0;
  assign T1028 = T1026[1'h0:1'h0];
  assign T1029 = T1026[1'h1:1'h1];
  assign T1030 = T1026[2'h2:2'h2];
  assign T1031 = T1038 ? creditConsReady_4_1 : T1032;
  assign T1032 = T1037 ? T1035 : T1033;
  assign T1033 = T1034 ? creditConsReady_1_1 : creditConsReady_0_1;
  assign T1034 = T1026[1'h0:1'h0];
  assign T1035 = T1036 ? creditConsReady_3_1 : creditConsReady_2_1;
  assign T1036 = T1026[1'h0:1'h0];
  assign T1037 = T1026[1'h1:1'h1];
  assign T1038 = T1026[2'h2:2'h2];
  assign T1039 = T3151;
  assign T3151 = R1002[1'h0:1'h0];
  assign T1040 = T1051 & T1041;
  assign T1041 = T1042 == 4'h4;
  assign T1042 = T1050 ? swAllocator_io_chosens_4 : T1043;
  assign T1043 = T1049 ? T1047 : T1044;
  assign T1044 = T1045 ? swAllocator_io_chosens_1 : swAllocator_io_chosens_0;
  assign T1045 = T1046[1'h0:1'h0];
  assign T1046 = R1015;
  assign T1047 = T1048 ? swAllocator_io_chosens_3 : swAllocator_io_chosens_2;
  assign T1048 = T1046[1'h0:1'h0];
  assign T1049 = T1046[1'h1:1'h1];
  assign T1050 = T1046[2'h2:2'h2];
  assign T1051 = T1059 ? swAllocator_io_requests_4_4_grant : T1052;
  assign T1052 = T1058 ? T1056 : T1053;
  assign T1053 = T1054 ? swAllocator_io_requests_1_4_grant : swAllocator_io_requests_0_4_grant;
  assign T1054 = T1055[1'h0:1'h0];
  assign T1055 = R1015;
  assign T1056 = T1057 ? swAllocator_io_requests_3_4_grant : swAllocator_io_requests_2_4_grant;
  assign T1057 = T1055[1'h0:1'h0];
  assign T1058 = T1055[1'h1:1'h1];
  assign T1059 = T1055[2'h2:2'h2];
  assign T1060 = RouterBuffer_4_io_deq_valid & T1061;
  assign T1061 = T1062;
  assign T1062 = T1067 ? T1065 : T1063;
  assign T1063 = T1064[6'h25:6'h25];
  assign T1064 = RouterBuffer_4_io_deq_bits_x[6'h36:1'h1];
  assign T1065 = T1066[4'he:4'he];
  assign T1066 = RouterBuffer_4_io_deq_bits_x[5'h1f:1'h1];
  assign T1067 = T1068 == 1'h1;
  assign T1068 = RouterBuffer_4_io_deq_bits_x[1'h0:1'h0];
  assign T3152 = reset ? 1'h0 : RouterBuffer_4_io_deq_valid;
  assign T1070 = T1071[2'h2:1'h0];
  assign T1071 = T1072[5'h1f:1'h1];
  assign T1072 = RouterRegFile_4_io_readData;
  assign T1073 = T1071[3'h4:2'h3];
  assign T1074 = T1071[3'h6:3'h5];
  assign T1075 = T1071[4'h8:3'h7];
  assign T1076 = T1071[4'hc:4'h9];
  assign T1077 = T1071[4'hd:4'hd];
  assign T1078 = T1071[4'he:4'he];
  assign T1079 = T1071[5'h1e:4'hf];
  assign T1080 = T1094 ? T1091 : T1081;
  assign T1081 = T1087 ? 1'h0 : T1082;
  assign T1082 = T1083 & T1021;
  assign T1083 = T1085 & T1084;
  assign T1084 = VCRouterStateManagement_4_io_currentState == 3'h4;
  assign T1085 = T1040 | T1086;
  assign T1086 = VCRouterStateManagement_4_io_currentState == 3'h4;
  assign T1087 = T1089 & T1088;
  assign T1088 = ~ RouterRegFile_4_io_readValid;
  assign T1089 = T1090 == 1'h1;
  assign T1090 = RouterBuffer_4_io_deq_bits_x[1'h0:1'h0];
  assign T1091 = T1092 & T1021;
  assign T1092 = T1085 & T1093;
  assign T1093 = 3'h3 <= VCRouterStateManagement_4_io_currentState;
  assign T1094 = T1098 & T1095;
  assign T1095 = T1096 & RouterRegFile_4_io_readValid;
  assign T1096 = T1097 == 1'h1;
  assign T1097 = RouterBuffer_4_io_deq_bits_x[1'h0:1'h0];
  assign T1098 = T1087 ^ 1'h1;
  assign T1099 = io_inChannels_2_flitValid & T114;
  assign T1100 = T1101 & RouterRegFile_4_io_readValid;
  assign T1101 = RouterRegFile_4_io_rvPipelineReg_0 ^ 1'h1;
  assign T1102 = T1104 & T1103;
  assign T1103 = VCRouterStateManagement_4_io_currentState == 3'h2;
  assign T1104 = RouterRegFile_4_io_rvPipelineReg_0 & vcAllocator_io_resources_4_valid;
  assign T1105 = T1107 & T1106;
  assign T1106 = VCRouterStateManagement_4_io_currentState == 3'h3;
  assign T1107 = RouterRegFile_4_io_rvPipelineReg_1 & T1040;
  assign T3153 = {24'h0, T1108};
  assign T1108 = T1109;
  assign T1109 = {T1113, T1110};
  assign T1110 = {T1112, T1111};
  assign T1111 = {CMeshDOR_4_io_outHeadFlit_destination_0, CMeshDOR_4_io_outHeadFlit_priorityLevel};
  assign T1112 = {CMeshDOR_4_io_outHeadFlit_destination_2, CMeshDOR_4_io_outHeadFlit_destination_1};
  assign T1113 = {T1115, T1114};
  assign T1114 = {CMeshDOR_4_io_outHeadFlit_vcPort, CMeshDOR_4_io_outHeadFlit_packetType};
  assign T1115 = {CMeshDOR_4_io_outHeadFlit_packetID, CMeshDOR_4_io_outHeadFlit_isTail};
  assign T1116 = T1118 & T1117;
  assign T1117 = VCRouterStateManagement_4_io_currentState == 3'h4;
  assign T1118 = T1119 & T1021;
  assign T1119 = T1085 & flitsAreTail_4;
  assign flitsAreTail_4 = T1120;
  assign T1120 = T1121 & RouterBuffer_4_io_deq_valid;
  assign T1121 = T1122;
  assign T1122 = T1127 ? T1125 : T1123;
  assign T1123 = T1124[6'h25:6'h25];
  assign T1124 = RouterBuffer_4_io_deq_bits_x[6'h36:1'h1];
  assign T1125 = T1126[4'he:4'he];
  assign T1126 = RouterBuffer_4_io_deq_bits_x[5'h1f:1'h1];
  assign T1127 = T1128 == 1'h1;
  assign T1128 = RouterBuffer_4_io_deq_bits_x[1'h0:1'h0];
  assign T1129 = T1130 ? T1099 : 1'h0;
  assign T1130 = T1131 == 1'h1;
  assign T1131 = io_inChannels_2_flit_x[1'h0:1'h0];
  assign T1132 = T1130 ? T1133 : 55'h0;
  assign T1133 = io_inChannels_2_flit_x;
  assign T1134 = T1094 ? T1140 : T1135;
  assign T1135 = T1087 ? 1'h0 : T1136;
  assign T1136 = T1137 & RouterBuffer_4_io_deq_valid;
  assign T1137 = T1138 & T1021;
  assign T1138 = T1085 & T1139;
  assign T1139 = VCRouterStateManagement_4_io_currentState == 3'h4;
  assign T1140 = T1141 & RouterBuffer_4_io_deq_valid;
  assign T1141 = T1142 & T1021;
  assign T1142 = T1085 & T1143;
  assign T1143 = 3'h3 <= VCRouterStateManagement_4_io_currentState;
  assign T1144 = T1145;
  assign T1145 = io_inChannels_1_flit_x;
  assign T3154 = R1146[1'h0:1'h0];
  assign T3155 = reset ? 55'h0 : T1147;
  assign T1147 = T1148 ? T3156 : R1146;
  assign T3156 = {51'h0, vcAllocator_io_chosens_3};
  assign T1148 = T1149 & vcAllocator_io_resources_3_valid;
  assign T1149 = VCRouterStateManagement_3_io_currentState == 3'h2;
  assign T1150 = T1151;
  assign T1151 = RouterBuffer_3_io_deq_bits_x;
  assign T1152 = T1164 | T1153;
  assign T1153 = T1154 == 2'h1;
  assign T1154 = T1163 ? VCRouterOutputStateManagement_4_io_currentState : T1155;
  assign T1155 = T1162 ? T1160 : T1156;
  assign T1156 = T1157 ? VCRouterOutputStateManagement_1_io_currentState : VCRouterOutputStateManagement_io_currentState;
  assign T1157 = T1158[1'h0:1'h0];
  assign T1158 = R1159;
  assign T3157 = reset ? 3'h0 : CMeshDOR_3_io_result;
  assign T1160 = T1161 ? VCRouterOutputStateManagement_3_io_currentState : VCRouterOutputStateManagement_2_io_currentState;
  assign T1161 = T1158[1'h0:1'h0];
  assign T1162 = T1158[1'h1:1'h1];
  assign T1163 = T1158[2'h2:2'h2];
  assign T1164 = T1154 == 2'h2;
  assign T1165 = T1183 ? T1175 : T1166;
  assign T1166 = T1174 ? creditConsReady_4_0 : T1167;
  assign T1167 = T1173 ? T1171 : T1168;
  assign T1168 = T1169 ? creditConsReady_1_0 : creditConsReady_0_0;
  assign T1169 = T1170[1'h0:1'h0];
  assign T1170 = R1159;
  assign T1171 = T1172 ? creditConsReady_3_0 : creditConsReady_2_0;
  assign T1172 = T1170[1'h0:1'h0];
  assign T1173 = T1170[1'h1:1'h1];
  assign T1174 = T1170[2'h2:2'h2];
  assign T1175 = T1182 ? creditConsReady_4_1 : T1176;
  assign T1176 = T1181 ? T1179 : T1177;
  assign T1177 = T1178 ? creditConsReady_1_1 : creditConsReady_0_1;
  assign T1178 = T1170[1'h0:1'h0];
  assign T1179 = T1180 ? creditConsReady_3_1 : creditConsReady_2_1;
  assign T1180 = T1170[1'h0:1'h0];
  assign T1181 = T1170[1'h1:1'h1];
  assign T1182 = T1170[2'h2:2'h2];
  assign T1183 = T3158;
  assign T3158 = R1146[1'h0:1'h0];
  assign T1184 = T1195 & T1185;
  assign T1185 = T1186 == 4'h3;
  assign T1186 = T1194 ? swAllocator_io_chosens_4 : T1187;
  assign T1187 = T1193 ? T1191 : T1188;
  assign T1188 = T1189 ? swAllocator_io_chosens_1 : swAllocator_io_chosens_0;
  assign T1189 = T1190[1'h0:1'h0];
  assign T1190 = R1159;
  assign T1191 = T1192 ? swAllocator_io_chosens_3 : swAllocator_io_chosens_2;
  assign T1192 = T1190[1'h0:1'h0];
  assign T1193 = T1190[1'h1:1'h1];
  assign T1194 = T1190[2'h2:2'h2];
  assign T1195 = T1203 ? swAllocator_io_requests_4_3_grant : T1196;
  assign T1196 = T1202 ? T1200 : T1197;
  assign T1197 = T1198 ? swAllocator_io_requests_1_3_grant : swAllocator_io_requests_0_3_grant;
  assign T1198 = T1199[1'h0:1'h0];
  assign T1199 = R1159;
  assign T1200 = T1201 ? swAllocator_io_requests_3_3_grant : swAllocator_io_requests_2_3_grant;
  assign T1201 = T1199[1'h0:1'h0];
  assign T1202 = T1199[1'h1:1'h1];
  assign T1203 = T1199[2'h2:2'h2];
  assign T1204 = RouterBuffer_3_io_deq_valid & T1205;
  assign T1205 = T1206;
  assign T1206 = T1211 ? T1209 : T1207;
  assign T1207 = T1208[6'h25:6'h25];
  assign T1208 = RouterBuffer_3_io_deq_bits_x[6'h36:1'h1];
  assign T1209 = T1210[4'he:4'he];
  assign T1210 = RouterBuffer_3_io_deq_bits_x[5'h1f:1'h1];
  assign T1211 = T1212 == 1'h1;
  assign T1212 = RouterBuffer_3_io_deq_bits_x[1'h0:1'h0];
  assign T3159 = reset ? 1'h0 : RouterBuffer_3_io_deq_valid;
  assign T1214 = T1215[2'h2:1'h0];
  assign T1215 = T1216[5'h1f:1'h1];
  assign T1216 = RouterRegFile_3_io_readData;
  assign T1217 = T1215[3'h4:2'h3];
  assign T1218 = T1215[3'h6:3'h5];
  assign T1219 = T1215[4'h8:3'h7];
  assign T1220 = T1215[4'hc:4'h9];
  assign T1221 = T1215[4'hd:4'hd];
  assign T1222 = T1215[4'he:4'he];
  assign T1223 = T1215[5'h1e:4'hf];
  assign T1224 = T1238 ? T1235 : T1225;
  assign T1225 = T1231 ? 1'h0 : T1226;
  assign T1226 = T1227 & T1165;
  assign T1227 = T1229 & T1228;
  assign T1228 = VCRouterStateManagement_3_io_currentState == 3'h4;
  assign T1229 = T1184 | T1230;
  assign T1230 = VCRouterStateManagement_3_io_currentState == 3'h4;
  assign T1231 = T1233 & T1232;
  assign T1232 = ~ RouterRegFile_3_io_readValid;
  assign T1233 = T1234 == 1'h1;
  assign T1234 = RouterBuffer_3_io_deq_bits_x[1'h0:1'h0];
  assign T1235 = T1236 & T1165;
  assign T1236 = T1229 & T1237;
  assign T1237 = 3'h3 <= VCRouterStateManagement_3_io_currentState;
  assign T1238 = T1242 & T1239;
  assign T1239 = T1240 & RouterRegFile_3_io_readValid;
  assign T1240 = T1241 == 1'h1;
  assign T1241 = RouterBuffer_3_io_deq_bits_x[1'h0:1'h0];
  assign T1242 = T1231 ^ 1'h1;
  assign T1243 = io_inChannels_1_flitValid & T136;
  assign T1244 = T1245 & RouterRegFile_3_io_readValid;
  assign T1245 = RouterRegFile_3_io_rvPipelineReg_0 ^ 1'h1;
  assign T1246 = T1248 & T1247;
  assign T1247 = VCRouterStateManagement_3_io_currentState == 3'h2;
  assign T1248 = RouterRegFile_3_io_rvPipelineReg_0 & vcAllocator_io_resources_3_valid;
  assign T1249 = T1251 & T1250;
  assign T1250 = VCRouterStateManagement_3_io_currentState == 3'h3;
  assign T1251 = RouterRegFile_3_io_rvPipelineReg_1 & T1184;
  assign T3160 = {24'h0, T1252};
  assign T1252 = T1253;
  assign T1253 = {T1257, T1254};
  assign T1254 = {T1256, T1255};
  assign T1255 = {CMeshDOR_3_io_outHeadFlit_destination_0, CMeshDOR_3_io_outHeadFlit_priorityLevel};
  assign T1256 = {CMeshDOR_3_io_outHeadFlit_destination_2, CMeshDOR_3_io_outHeadFlit_destination_1};
  assign T1257 = {T1259, T1258};
  assign T1258 = {CMeshDOR_3_io_outHeadFlit_vcPort, CMeshDOR_3_io_outHeadFlit_packetType};
  assign T1259 = {CMeshDOR_3_io_outHeadFlit_packetID, CMeshDOR_3_io_outHeadFlit_isTail};
  assign T1260 = T1262 & T1261;
  assign T1261 = VCRouterStateManagement_3_io_currentState == 3'h4;
  assign T1262 = T1263 & T1165;
  assign T1263 = T1229 & flitsAreTail_3;
  assign flitsAreTail_3 = T1264;
  assign T1264 = T1265 & RouterBuffer_3_io_deq_valid;
  assign T1265 = T1266;
  assign T1266 = T1271 ? T1269 : T1267;
  assign T1267 = T1268[6'h25:6'h25];
  assign T1268 = RouterBuffer_3_io_deq_bits_x[6'h36:1'h1];
  assign T1269 = T1270[4'he:4'he];
  assign T1270 = RouterBuffer_3_io_deq_bits_x[5'h1f:1'h1];
  assign T1271 = T1272 == 1'h1;
  assign T1272 = RouterBuffer_3_io_deq_bits_x[1'h0:1'h0];
  assign T1273 = T1274 ? T1243 : 1'h0;
  assign T1274 = T1275 == 1'h1;
  assign T1275 = io_inChannels_1_flit_x[1'h0:1'h0];
  assign T1276 = T1274 ? T1277 : 55'h0;
  assign T1277 = io_inChannels_1_flit_x;
  assign T1278 = T1238 ? T1284 : T1279;
  assign T1279 = T1231 ? 1'h0 : T1280;
  assign T1280 = T1281 & RouterBuffer_3_io_deq_valid;
  assign T1281 = T1282 & T1165;
  assign T1282 = T1229 & T1283;
  assign T1283 = VCRouterStateManagement_3_io_currentState == 3'h4;
  assign T1284 = T1285 & RouterBuffer_3_io_deq_valid;
  assign T1285 = T1286 & T1165;
  assign T1286 = T1229 & T1287;
  assign T1287 = 3'h3 <= VCRouterStateManagement_3_io_currentState;
  assign T1288 = T1289;
  assign T1289 = io_inChannels_1_flit_x;
  assign T3161 = R1290[1'h0:1'h0];
  assign T3162 = reset ? 55'h0 : T1291;
  assign T1291 = T1292 ? T3163 : R1290;
  assign T3163 = {51'h0, vcAllocator_io_chosens_2};
  assign T1292 = T1293 & vcAllocator_io_resources_2_valid;
  assign T1293 = VCRouterStateManagement_2_io_currentState == 3'h2;
  assign T1294 = T1295;
  assign T1295 = RouterBuffer_2_io_deq_bits_x;
  assign T1296 = T1308 | T1297;
  assign T1297 = T1298 == 2'h1;
  assign T1298 = T1307 ? VCRouterOutputStateManagement_4_io_currentState : T1299;
  assign T1299 = T1306 ? T1304 : T1300;
  assign T1300 = T1301 ? VCRouterOutputStateManagement_1_io_currentState : VCRouterOutputStateManagement_io_currentState;
  assign T1301 = T1302[1'h0:1'h0];
  assign T1302 = R1303;
  assign T3164 = reset ? 3'h0 : CMeshDOR_2_io_result;
  assign T1304 = T1305 ? VCRouterOutputStateManagement_3_io_currentState : VCRouterOutputStateManagement_2_io_currentState;
  assign T1305 = T1302[1'h0:1'h0];
  assign T1306 = T1302[1'h1:1'h1];
  assign T1307 = T1302[2'h2:2'h2];
  assign T1308 = T1298 == 2'h2;
  assign T1309 = T1327 ? T1319 : T1310;
  assign T1310 = T1318 ? creditConsReady_4_0 : T1311;
  assign T1311 = T1317 ? T1315 : T1312;
  assign T1312 = T1313 ? creditConsReady_1_0 : creditConsReady_0_0;
  assign T1313 = T1314[1'h0:1'h0];
  assign T1314 = R1303;
  assign T1315 = T1316 ? creditConsReady_3_0 : creditConsReady_2_0;
  assign T1316 = T1314[1'h0:1'h0];
  assign T1317 = T1314[1'h1:1'h1];
  assign T1318 = T1314[2'h2:2'h2];
  assign T1319 = T1326 ? creditConsReady_4_1 : T1320;
  assign T1320 = T1325 ? T1323 : T1321;
  assign T1321 = T1322 ? creditConsReady_1_1 : creditConsReady_0_1;
  assign T1322 = T1314[1'h0:1'h0];
  assign T1323 = T1324 ? creditConsReady_3_1 : creditConsReady_2_1;
  assign T1324 = T1314[1'h0:1'h0];
  assign T1325 = T1314[1'h1:1'h1];
  assign T1326 = T1314[2'h2:2'h2];
  assign T1327 = T3165;
  assign T3165 = R1290[1'h0:1'h0];
  assign T1328 = T1339 & T1329;
  assign T1329 = T1330 == 4'h2;
  assign T1330 = T1338 ? swAllocator_io_chosens_4 : T1331;
  assign T1331 = T1337 ? T1335 : T1332;
  assign T1332 = T1333 ? swAllocator_io_chosens_1 : swAllocator_io_chosens_0;
  assign T1333 = T1334[1'h0:1'h0];
  assign T1334 = R1303;
  assign T1335 = T1336 ? swAllocator_io_chosens_3 : swAllocator_io_chosens_2;
  assign T1336 = T1334[1'h0:1'h0];
  assign T1337 = T1334[1'h1:1'h1];
  assign T1338 = T1334[2'h2:2'h2];
  assign T1339 = T1347 ? swAllocator_io_requests_4_2_grant : T1340;
  assign T1340 = T1346 ? T1344 : T1341;
  assign T1341 = T1342 ? swAllocator_io_requests_1_2_grant : swAllocator_io_requests_0_2_grant;
  assign T1342 = T1343[1'h0:1'h0];
  assign T1343 = R1303;
  assign T1344 = T1345 ? swAllocator_io_requests_3_2_grant : swAllocator_io_requests_2_2_grant;
  assign T1345 = T1343[1'h0:1'h0];
  assign T1346 = T1343[1'h1:1'h1];
  assign T1347 = T1343[2'h2:2'h2];
  assign T1348 = RouterBuffer_2_io_deq_valid & T1349;
  assign T1349 = T1350;
  assign T1350 = T1355 ? T1353 : T1351;
  assign T1351 = T1352[6'h25:6'h25];
  assign T1352 = RouterBuffer_2_io_deq_bits_x[6'h36:1'h1];
  assign T1353 = T1354[4'he:4'he];
  assign T1354 = RouterBuffer_2_io_deq_bits_x[5'h1f:1'h1];
  assign T1355 = T1356 == 1'h1;
  assign T1356 = RouterBuffer_2_io_deq_bits_x[1'h0:1'h0];
  assign T3166 = reset ? 1'h0 : RouterBuffer_2_io_deq_valid;
  assign T1358 = T1359[2'h2:1'h0];
  assign T1359 = T1360[5'h1f:1'h1];
  assign T1360 = RouterRegFile_2_io_readData;
  assign T1361 = T1359[3'h4:2'h3];
  assign T1362 = T1359[3'h6:3'h5];
  assign T1363 = T1359[4'h8:3'h7];
  assign T1364 = T1359[4'hc:4'h9];
  assign T1365 = T1359[4'hd:4'hd];
  assign T1366 = T1359[4'he:4'he];
  assign T1367 = T1359[5'h1e:4'hf];
  assign T1368 = T1382 ? T1379 : T1369;
  assign T1369 = T1375 ? 1'h0 : T1370;
  assign T1370 = T1371 & T1309;
  assign T1371 = T1373 & T1372;
  assign T1372 = VCRouterStateManagement_2_io_currentState == 3'h4;
  assign T1373 = T1328 | T1374;
  assign T1374 = VCRouterStateManagement_2_io_currentState == 3'h4;
  assign T1375 = T1377 & T1376;
  assign T1376 = ~ RouterRegFile_2_io_readValid;
  assign T1377 = T1378 == 1'h1;
  assign T1378 = RouterBuffer_2_io_deq_bits_x[1'h0:1'h0];
  assign T1379 = T1380 & T1309;
  assign T1380 = T1373 & T1381;
  assign T1381 = 3'h3 <= VCRouterStateManagement_2_io_currentState;
  assign T1382 = T1386 & T1383;
  assign T1383 = T1384 & RouterRegFile_2_io_readValid;
  assign T1384 = T1385 == 1'h1;
  assign T1385 = RouterBuffer_2_io_deq_bits_x[1'h0:1'h0];
  assign T1386 = T1375 ^ 1'h1;
  assign T1387 = io_inChannels_1_flitValid & T158;
  assign T1388 = T1389 & RouterRegFile_2_io_readValid;
  assign T1389 = RouterRegFile_2_io_rvPipelineReg_0 ^ 1'h1;
  assign T1390 = T1392 & T1391;
  assign T1391 = VCRouterStateManagement_2_io_currentState == 3'h2;
  assign T1392 = RouterRegFile_2_io_rvPipelineReg_0 & vcAllocator_io_resources_2_valid;
  assign T1393 = T1395 & T1394;
  assign T1394 = VCRouterStateManagement_2_io_currentState == 3'h3;
  assign T1395 = RouterRegFile_2_io_rvPipelineReg_1 & T1328;
  assign T3167 = {24'h0, T1396};
  assign T1396 = T1397;
  assign T1397 = {T1401, T1398};
  assign T1398 = {T1400, T1399};
  assign T1399 = {CMeshDOR_2_io_outHeadFlit_destination_0, CMeshDOR_2_io_outHeadFlit_priorityLevel};
  assign T1400 = {CMeshDOR_2_io_outHeadFlit_destination_2, CMeshDOR_2_io_outHeadFlit_destination_1};
  assign T1401 = {T1403, T1402};
  assign T1402 = {CMeshDOR_2_io_outHeadFlit_vcPort, CMeshDOR_2_io_outHeadFlit_packetType};
  assign T1403 = {CMeshDOR_2_io_outHeadFlit_packetID, CMeshDOR_2_io_outHeadFlit_isTail};
  assign T1404 = T1406 & T1405;
  assign T1405 = VCRouterStateManagement_2_io_currentState == 3'h4;
  assign T1406 = T1407 & T1309;
  assign T1407 = T1373 & flitsAreTail_2;
  assign flitsAreTail_2 = T1408;
  assign T1408 = T1409 & RouterBuffer_2_io_deq_valid;
  assign T1409 = T1410;
  assign T1410 = T1415 ? T1413 : T1411;
  assign T1411 = T1412[6'h25:6'h25];
  assign T1412 = RouterBuffer_2_io_deq_bits_x[6'h36:1'h1];
  assign T1413 = T1414[4'he:4'he];
  assign T1414 = RouterBuffer_2_io_deq_bits_x[5'h1f:1'h1];
  assign T1415 = T1416 == 1'h1;
  assign T1416 = RouterBuffer_2_io_deq_bits_x[1'h0:1'h0];
  assign T1417 = T1418 ? T1387 : 1'h0;
  assign T1418 = T1419 == 1'h1;
  assign T1419 = io_inChannels_1_flit_x[1'h0:1'h0];
  assign T1420 = T1418 ? T1421 : 55'h0;
  assign T1421 = io_inChannels_1_flit_x;
  assign T1422 = T1382 ? T1428 : T1423;
  assign T1423 = T1375 ? 1'h0 : T1424;
  assign T1424 = T1425 & RouterBuffer_2_io_deq_valid;
  assign T1425 = T1426 & T1309;
  assign T1426 = T1373 & T1427;
  assign T1427 = VCRouterStateManagement_2_io_currentState == 3'h4;
  assign T1428 = T1429 & RouterBuffer_2_io_deq_valid;
  assign T1429 = T1430 & T1309;
  assign T1430 = T1373 & T1431;
  assign T1431 = 3'h3 <= VCRouterStateManagement_2_io_currentState;
  assign T1432 = T1433;
  assign T1433 = io_inChannels_0_flit_x;
  assign T3168 = R1434[1'h0:1'h0];
  assign T3169 = reset ? 55'h0 : T1435;
  assign T1435 = T1436 ? T3170 : R1434;
  assign T3170 = {51'h0, vcAllocator_io_chosens_1};
  assign T1436 = T1437 & vcAllocator_io_resources_1_valid;
  assign T1437 = VCRouterStateManagement_1_io_currentState == 3'h2;
  assign T1438 = T1439;
  assign T1439 = RouterBuffer_1_io_deq_bits_x;
  assign T1440 = T1452 | T1441;
  assign T1441 = T1442 == 2'h1;
  assign T1442 = T1451 ? VCRouterOutputStateManagement_4_io_currentState : T1443;
  assign T1443 = T1450 ? T1448 : T1444;
  assign T1444 = T1445 ? VCRouterOutputStateManagement_1_io_currentState : VCRouterOutputStateManagement_io_currentState;
  assign T1445 = T1446[1'h0:1'h0];
  assign T1446 = R1447;
  assign T3171 = reset ? 3'h0 : CMeshDOR_1_io_result;
  assign T1448 = T1449 ? VCRouterOutputStateManagement_3_io_currentState : VCRouterOutputStateManagement_2_io_currentState;
  assign T1449 = T1446[1'h0:1'h0];
  assign T1450 = T1446[1'h1:1'h1];
  assign T1451 = T1446[2'h2:2'h2];
  assign T1452 = T1442 == 2'h2;
  assign T1453 = T1471 ? T1463 : T1454;
  assign T1454 = T1462 ? creditConsReady_4_0 : T1455;
  assign T1455 = T1461 ? T1459 : T1456;
  assign T1456 = T1457 ? creditConsReady_1_0 : creditConsReady_0_0;
  assign T1457 = T1458[1'h0:1'h0];
  assign T1458 = R1447;
  assign T1459 = T1460 ? creditConsReady_3_0 : creditConsReady_2_0;
  assign T1460 = T1458[1'h0:1'h0];
  assign T1461 = T1458[1'h1:1'h1];
  assign T1462 = T1458[2'h2:2'h2];
  assign T1463 = T1470 ? creditConsReady_4_1 : T1464;
  assign T1464 = T1469 ? T1467 : T1465;
  assign T1465 = T1466 ? creditConsReady_1_1 : creditConsReady_0_1;
  assign T1466 = T1458[1'h0:1'h0];
  assign T1467 = T1468 ? creditConsReady_3_1 : creditConsReady_2_1;
  assign T1468 = T1458[1'h0:1'h0];
  assign T1469 = T1458[1'h1:1'h1];
  assign T1470 = T1458[2'h2:2'h2];
  assign T1471 = T3172;
  assign T3172 = R1434[1'h0:1'h0];
  assign T1472 = T1483 & T1473;
  assign T1473 = T1474 == 4'h1;
  assign T1474 = T1482 ? swAllocator_io_chosens_4 : T1475;
  assign T1475 = T1481 ? T1479 : T1476;
  assign T1476 = T1477 ? swAllocator_io_chosens_1 : swAllocator_io_chosens_0;
  assign T1477 = T1478[1'h0:1'h0];
  assign T1478 = R1447;
  assign T1479 = T1480 ? swAllocator_io_chosens_3 : swAllocator_io_chosens_2;
  assign T1480 = T1478[1'h0:1'h0];
  assign T1481 = T1478[1'h1:1'h1];
  assign T1482 = T1478[2'h2:2'h2];
  assign T1483 = T1491 ? swAllocator_io_requests_4_1_grant : T1484;
  assign T1484 = T1490 ? T1488 : T1485;
  assign T1485 = T1486 ? swAllocator_io_requests_1_1_grant : swAllocator_io_requests_0_1_grant;
  assign T1486 = T1487[1'h0:1'h0];
  assign T1487 = R1447;
  assign T1488 = T1489 ? swAllocator_io_requests_3_1_grant : swAllocator_io_requests_2_1_grant;
  assign T1489 = T1487[1'h0:1'h0];
  assign T1490 = T1487[1'h1:1'h1];
  assign T1491 = T1487[2'h2:2'h2];
  assign T1492 = RouterBuffer_1_io_deq_valid & T1493;
  assign T1493 = T1494;
  assign T1494 = T1499 ? T1497 : T1495;
  assign T1495 = T1496[6'h25:6'h25];
  assign T1496 = RouterBuffer_1_io_deq_bits_x[6'h36:1'h1];
  assign T1497 = T1498[4'he:4'he];
  assign T1498 = RouterBuffer_1_io_deq_bits_x[5'h1f:1'h1];
  assign T1499 = T1500 == 1'h1;
  assign T1500 = RouterBuffer_1_io_deq_bits_x[1'h0:1'h0];
  assign T3173 = reset ? 1'h0 : RouterBuffer_1_io_deq_valid;
  assign T1502 = T1503[2'h2:1'h0];
  assign T1503 = T1504[5'h1f:1'h1];
  assign T1504 = RouterRegFile_1_io_readData;
  assign T1505 = T1503[3'h4:2'h3];
  assign T1506 = T1503[3'h6:3'h5];
  assign T1507 = T1503[4'h8:3'h7];
  assign T1508 = T1503[4'hc:4'h9];
  assign T1509 = T1503[4'hd:4'hd];
  assign T1510 = T1503[4'he:4'he];
  assign T1511 = T1503[5'h1e:4'hf];
  assign T1512 = T1526 ? T1523 : T1513;
  assign T1513 = T1519 ? 1'h0 : T1514;
  assign T1514 = T1515 & T1453;
  assign T1515 = T1517 & T1516;
  assign T1516 = VCRouterStateManagement_1_io_currentState == 3'h4;
  assign T1517 = T1472 | T1518;
  assign T1518 = VCRouterStateManagement_1_io_currentState == 3'h4;
  assign T1519 = T1521 & T1520;
  assign T1520 = ~ RouterRegFile_1_io_readValid;
  assign T1521 = T1522 == 1'h1;
  assign T1522 = RouterBuffer_1_io_deq_bits_x[1'h0:1'h0];
  assign T1523 = T1524 & T1453;
  assign T1524 = T1517 & T1525;
  assign T1525 = 3'h3 <= VCRouterStateManagement_1_io_currentState;
  assign T1526 = T1530 & T1527;
  assign T1527 = T1528 & RouterRegFile_1_io_readValid;
  assign T1528 = T1529 == 1'h1;
  assign T1529 = RouterBuffer_1_io_deq_bits_x[1'h0:1'h0];
  assign T1530 = T1519 ^ 1'h1;
  assign T1531 = io_inChannels_0_flitValid & T180;
  assign T1532 = T1533 & RouterRegFile_1_io_readValid;
  assign T1533 = RouterRegFile_1_io_rvPipelineReg_0 ^ 1'h1;
  assign T1534 = T1536 & T1535;
  assign T1535 = VCRouterStateManagement_1_io_currentState == 3'h2;
  assign T1536 = RouterRegFile_1_io_rvPipelineReg_0 & vcAllocator_io_resources_1_valid;
  assign T1537 = T1539 & T1538;
  assign T1538 = VCRouterStateManagement_1_io_currentState == 3'h3;
  assign T1539 = RouterRegFile_1_io_rvPipelineReg_1 & T1472;
  assign T3174 = {24'h0, T1540};
  assign T1540 = T1541;
  assign T1541 = {T1545, T1542};
  assign T1542 = {T1544, T1543};
  assign T1543 = {CMeshDOR_1_io_outHeadFlit_destination_0, CMeshDOR_1_io_outHeadFlit_priorityLevel};
  assign T1544 = {CMeshDOR_1_io_outHeadFlit_destination_2, CMeshDOR_1_io_outHeadFlit_destination_1};
  assign T1545 = {T1547, T1546};
  assign T1546 = {CMeshDOR_1_io_outHeadFlit_vcPort, CMeshDOR_1_io_outHeadFlit_packetType};
  assign T1547 = {CMeshDOR_1_io_outHeadFlit_packetID, CMeshDOR_1_io_outHeadFlit_isTail};
  assign T1548 = T1550 & T1549;
  assign T1549 = VCRouterStateManagement_1_io_currentState == 3'h4;
  assign T1550 = T1551 & T1453;
  assign T1551 = T1517 & flitsAreTail_1;
  assign flitsAreTail_1 = T1552;
  assign T1552 = T1553 & RouterBuffer_1_io_deq_valid;
  assign T1553 = T1554;
  assign T1554 = T1559 ? T1557 : T1555;
  assign T1555 = T1556[6'h25:6'h25];
  assign T1556 = RouterBuffer_1_io_deq_bits_x[6'h36:1'h1];
  assign T1557 = T1558[4'he:4'he];
  assign T1558 = RouterBuffer_1_io_deq_bits_x[5'h1f:1'h1];
  assign T1559 = T1560 == 1'h1;
  assign T1560 = RouterBuffer_1_io_deq_bits_x[1'h0:1'h0];
  assign T1561 = T1562 ? T1531 : 1'h0;
  assign T1562 = T1563 == 1'h1;
  assign T1563 = io_inChannels_0_flit_x[1'h0:1'h0];
  assign T1564 = T1562 ? T1565 : 55'h0;
  assign T1565 = io_inChannels_0_flit_x;
  assign T1566 = T1526 ? T1572 : T1567;
  assign T1567 = T1519 ? 1'h0 : T1568;
  assign T1568 = T1569 & RouterBuffer_1_io_deq_valid;
  assign T1569 = T1570 & T1453;
  assign T1570 = T1517 & T1571;
  assign T1571 = VCRouterStateManagement_1_io_currentState == 3'h4;
  assign T1572 = T1573 & RouterBuffer_1_io_deq_valid;
  assign T1573 = T1574 & T1453;
  assign T1574 = T1517 & T1575;
  assign T1575 = 3'h3 <= VCRouterStateManagement_1_io_currentState;
  assign T1576 = T1577;
  assign T1577 = io_inChannels_0_flit_x;
  assign T3175 = R1578[1'h0:1'h0];
  assign T3176 = reset ? 55'h0 : T1579;
  assign T1579 = T1580 ? T3177 : R1578;
  assign T3177 = {51'h0, vcAllocator_io_chosens_0};
  assign T1580 = T1581 & vcAllocator_io_resources_0_valid;
  assign T1581 = VCRouterStateManagement_io_currentState == 3'h2;
  assign T1582 = T1583;
  assign T1583 = RouterBuffer_io_deq_bits_x;
  assign T1584 = T1596 | T1585;
  assign T1585 = T1586 == 2'h1;
  assign T1586 = T1595 ? VCRouterOutputStateManagement_4_io_currentState : T1587;
  assign T1587 = T1594 ? T1592 : T1588;
  assign T1588 = T1589 ? VCRouterOutputStateManagement_1_io_currentState : VCRouterOutputStateManagement_io_currentState;
  assign T1589 = T1590[1'h0:1'h0];
  assign T1590 = R1591;
  assign T3178 = reset ? 3'h0 : CMeshDOR_io_result;
  assign T1592 = T1593 ? VCRouterOutputStateManagement_3_io_currentState : VCRouterOutputStateManagement_2_io_currentState;
  assign T1593 = T1590[1'h0:1'h0];
  assign T1594 = T1590[1'h1:1'h1];
  assign T1595 = T1590[2'h2:2'h2];
  assign T1596 = T1586 == 2'h2;
  assign T1597 = T1615 ? T1607 : T1598;
  assign T1598 = T1606 ? creditConsReady_4_0 : T1599;
  assign T1599 = T1605 ? T1603 : T1600;
  assign T1600 = T1601 ? creditConsReady_1_0 : creditConsReady_0_0;
  assign T1601 = T1602[1'h0:1'h0];
  assign T1602 = R1591;
  assign T1603 = T1604 ? creditConsReady_3_0 : creditConsReady_2_0;
  assign T1604 = T1602[1'h0:1'h0];
  assign T1605 = T1602[1'h1:1'h1];
  assign T1606 = T1602[2'h2:2'h2];
  assign T1607 = T1614 ? creditConsReady_4_1 : T1608;
  assign T1608 = T1613 ? T1611 : T1609;
  assign T1609 = T1610 ? creditConsReady_1_1 : creditConsReady_0_1;
  assign T1610 = T1602[1'h0:1'h0];
  assign T1611 = T1612 ? creditConsReady_3_1 : creditConsReady_2_1;
  assign T1612 = T1602[1'h0:1'h0];
  assign T1613 = T1602[1'h1:1'h1];
  assign T1614 = T1602[2'h2:2'h2];
  assign T1615 = T3179;
  assign T3179 = R1578[1'h0:1'h0];
  assign T1616 = T1627 & T1617;
  assign T1617 = T1618 == 4'h0;
  assign T1618 = T1626 ? swAllocator_io_chosens_4 : T1619;
  assign T1619 = T1625 ? T1623 : T1620;
  assign T1620 = T1621 ? swAllocator_io_chosens_1 : swAllocator_io_chosens_0;
  assign T1621 = T1622[1'h0:1'h0];
  assign T1622 = R1591;
  assign T1623 = T1624 ? swAllocator_io_chosens_3 : swAllocator_io_chosens_2;
  assign T1624 = T1622[1'h0:1'h0];
  assign T1625 = T1622[1'h1:1'h1];
  assign T1626 = T1622[2'h2:2'h2];
  assign T1627 = T1635 ? swAllocator_io_requests_4_0_grant : T1628;
  assign T1628 = T1634 ? T1632 : T1629;
  assign T1629 = T1630 ? swAllocator_io_requests_1_0_grant : swAllocator_io_requests_0_0_grant;
  assign T1630 = T1631[1'h0:1'h0];
  assign T1631 = R1591;
  assign T1632 = T1633 ? swAllocator_io_requests_3_0_grant : swAllocator_io_requests_2_0_grant;
  assign T1633 = T1631[1'h0:1'h0];
  assign T1634 = T1631[1'h1:1'h1];
  assign T1635 = T1631[2'h2:2'h2];
  assign T1636 = RouterBuffer_io_deq_valid & T1637;
  assign T1637 = T1638;
  assign T1638 = T1643 ? T1641 : T1639;
  assign T1639 = T1640[6'h25:6'h25];
  assign T1640 = RouterBuffer_io_deq_bits_x[6'h36:1'h1];
  assign T1641 = T1642[4'he:4'he];
  assign T1642 = RouterBuffer_io_deq_bits_x[5'h1f:1'h1];
  assign T1643 = T1644 == 1'h1;
  assign T1644 = RouterBuffer_io_deq_bits_x[1'h0:1'h0];
  assign T3180 = reset ? 1'h0 : RouterBuffer_io_deq_valid;
  assign T1646 = T1647[2'h2:1'h0];
  assign T1647 = T1648[5'h1f:1'h1];
  assign T1648 = RouterRegFile_io_readData;
  assign T1649 = T1647[3'h4:2'h3];
  assign T1650 = T1647[3'h6:3'h5];
  assign T1651 = T1647[4'h8:3'h7];
  assign T1652 = T1647[4'hc:4'h9];
  assign T1653 = T1647[4'hd:4'hd];
  assign T1654 = T1647[4'he:4'he];
  assign T1655 = T1647[5'h1e:4'hf];
  assign T1656 = T1670 ? T1667 : T1657;
  assign T1657 = T1663 ? 1'h0 : T1658;
  assign T1658 = T1659 & T1597;
  assign T1659 = T1661 & T1660;
  assign T1660 = VCRouterStateManagement_io_currentState == 3'h4;
  assign T1661 = T1616 | T1662;
  assign T1662 = VCRouterStateManagement_io_currentState == 3'h4;
  assign T1663 = T1665 & T1664;
  assign T1664 = ~ RouterRegFile_io_readValid;
  assign T1665 = T1666 == 1'h1;
  assign T1666 = RouterBuffer_io_deq_bits_x[1'h0:1'h0];
  assign T1667 = T1668 & T1597;
  assign T1668 = T1661 & T1669;
  assign T1669 = 3'h3 <= VCRouterStateManagement_io_currentState;
  assign T1670 = T1674 & T1671;
  assign T1671 = T1672 & RouterRegFile_io_readValid;
  assign T1672 = T1673 == 1'h1;
  assign T1673 = RouterBuffer_io_deq_bits_x[1'h0:1'h0];
  assign T1674 = T1663 ^ 1'h1;
  assign T1675 = io_inChannels_0_flitValid & T202;
  assign T1676 = T1677 & RouterRegFile_io_readValid;
  assign T1677 = RouterRegFile_io_rvPipelineReg_0 ^ 1'h1;
  assign T1678 = T1680 & T1679;
  assign T1679 = VCRouterStateManagement_io_currentState == 3'h2;
  assign T1680 = RouterRegFile_io_rvPipelineReg_0 & vcAllocator_io_resources_0_valid;
  assign T1681 = T1683 & T1682;
  assign T1682 = VCRouterStateManagement_io_currentState == 3'h3;
  assign T1683 = RouterRegFile_io_rvPipelineReg_1 & T1616;
  assign T3181 = {24'h0, T1684};
  assign T1684 = T1685;
  assign T1685 = {T1689, T1686};
  assign T1686 = {T1688, T1687};
  assign T1687 = {CMeshDOR_io_outHeadFlit_destination_0, CMeshDOR_io_outHeadFlit_priorityLevel};
  assign T1688 = {CMeshDOR_io_outHeadFlit_destination_2, CMeshDOR_io_outHeadFlit_destination_1};
  assign T1689 = {T1691, T1690};
  assign T1690 = {CMeshDOR_io_outHeadFlit_vcPort, CMeshDOR_io_outHeadFlit_packetType};
  assign T1691 = {CMeshDOR_io_outHeadFlit_packetID, CMeshDOR_io_outHeadFlit_isTail};
  assign T1692 = T1694 & T1693;
  assign T1693 = VCRouterStateManagement_io_currentState == 3'h4;
  assign T1694 = T1695 & T1597;
  assign T1695 = T1661 & flitsAreTail_0;
  assign flitsAreTail_0 = T1696;
  assign T1696 = T1697 & RouterBuffer_io_deq_valid;
  assign T1697 = T1698;
  assign T1698 = T1703 ? T1701 : T1699;
  assign T1699 = T1700[6'h25:6'h25];
  assign T1700 = RouterBuffer_io_deq_bits_x[6'h36:1'h1];
  assign T1701 = T1702[4'he:4'he];
  assign T1702 = RouterBuffer_io_deq_bits_x[5'h1f:1'h1];
  assign T1703 = T1704 == 1'h1;
  assign T1704 = RouterBuffer_io_deq_bits_x[1'h0:1'h0];
  assign T1705 = T1706 ? T1675 : 1'h0;
  assign T1706 = T1707 == 1'h1;
  assign T1707 = io_inChannels_0_flit_x[1'h0:1'h0];
  assign T1708 = T1706 ? T1709 : 55'h0;
  assign T1709 = io_inChannels_0_flit_x;
  assign T1710 = T1670 ? T1716 : T1711;
  assign T1711 = T1663 ? 1'h0 : T1712;
  assign T1712 = T1713 & RouterBuffer_io_deq_valid;
  assign T1713 = T1714 & T1597;
  assign T1714 = T1661 & T1715;
  assign T1715 = VCRouterStateManagement_io_currentState == 3'h4;
  assign T1716 = T1717 & RouterBuffer_io_deq_valid;
  assign T1717 = T1718 & T1597;
  assign T1718 = T1661 & T1719;
  assign T1719 = 3'h3 <= VCRouterStateManagement_io_currentState;
  assign T1720 = T1721 ? CreditCon_9_io_outCredit : CreditCon_8_io_outCredit;
  assign T1721 = T222;
  assign T1722 = T1723 != 10'h0;
  assign T1723 = T1724;
  assign T1724 = {T1814, T1725};
  assign T1725 = {T1779, T1726};
  assign T1726 = {readyToXmit_2_4, T1727};
  assign T1727 = {readyToXmit_1_4, readyToXmit_0_4};
  assign readyToXmit_0_4 = T1728;
  assign T1728 = T1742 ? T1738 : T1729;
  assign T1729 = T1734 ? T1730 : 1'h0;
  assign T1730 = T1731 & RouterBuffer_io_deq_valid;
  assign T1731 = T1732 & T1597;
  assign T1732 = T1661 & T1733;
  assign T1733 = 3'h3 <= VCRouterStateManagement_io_currentState;
  assign T1734 = T1670 & T1735;
  assign T1735 = T1736[3'h4:3'h4];
  assign T1736 = 1'h1 << T1737;
  assign T1737 = R1591;
  assign T1738 = T1739 & RouterBuffer_io_deq_valid;
  assign T1739 = T1740 & T1597;
  assign T1740 = T1661 & T1741;
  assign T1741 = VCRouterStateManagement_io_currentState == 3'h4;
  assign T1742 = T1743 & T1735;
  assign T1743 = T1744 ^ 1'h1;
  assign T1744 = T1663 | T1671;
  assign readyToXmit_1_4 = T1745;
  assign T1745 = T1759 ? T1755 : T1746;
  assign T1746 = T1751 ? T1747 : 1'h0;
  assign T1747 = T1748 & RouterBuffer_1_io_deq_valid;
  assign T1748 = T1749 & T1453;
  assign T1749 = T1517 & T1750;
  assign T1750 = 3'h3 <= VCRouterStateManagement_1_io_currentState;
  assign T1751 = T1526 & T1752;
  assign T1752 = T1753[3'h4:3'h4];
  assign T1753 = 1'h1 << T1754;
  assign T1754 = R1447;
  assign T1755 = T1756 & RouterBuffer_1_io_deq_valid;
  assign T1756 = T1757 & T1453;
  assign T1757 = T1517 & T1758;
  assign T1758 = VCRouterStateManagement_1_io_currentState == 3'h4;
  assign T1759 = T1760 & T1752;
  assign T1760 = T1761 ^ 1'h1;
  assign T1761 = T1519 | T1527;
  assign readyToXmit_2_4 = T1762;
  assign T1762 = T1776 ? T1772 : T1763;
  assign T1763 = T1768 ? T1764 : 1'h0;
  assign T1764 = T1765 & RouterBuffer_2_io_deq_valid;
  assign T1765 = T1766 & T1309;
  assign T1766 = T1373 & T1767;
  assign T1767 = 3'h3 <= VCRouterStateManagement_2_io_currentState;
  assign T1768 = T1382 & T1769;
  assign T1769 = T1770[3'h4:3'h4];
  assign T1770 = 1'h1 << T1771;
  assign T1771 = R1303;
  assign T1772 = T1773 & RouterBuffer_2_io_deq_valid;
  assign T1773 = T1774 & T1309;
  assign T1774 = T1373 & T1775;
  assign T1775 = VCRouterStateManagement_2_io_currentState == 3'h4;
  assign T1776 = T1777 & T1769;
  assign T1777 = T1778 ^ 1'h1;
  assign T1778 = T1375 | T1383;
  assign T1779 = {readyToXmit_4_4, readyToXmit_3_4};
  assign readyToXmit_3_4 = T1780;
  assign T1780 = T1794 ? T1790 : T1781;
  assign T1781 = T1786 ? T1782 : 1'h0;
  assign T1782 = T1783 & RouterBuffer_3_io_deq_valid;
  assign T1783 = T1784 & T1165;
  assign T1784 = T1229 & T1785;
  assign T1785 = 3'h3 <= VCRouterStateManagement_3_io_currentState;
  assign T1786 = T1238 & T1787;
  assign T1787 = T1788[3'h4:3'h4];
  assign T1788 = 1'h1 << T1789;
  assign T1789 = R1159;
  assign T1790 = T1791 & RouterBuffer_3_io_deq_valid;
  assign T1791 = T1792 & T1165;
  assign T1792 = T1229 & T1793;
  assign T1793 = VCRouterStateManagement_3_io_currentState == 3'h4;
  assign T1794 = T1795 & T1787;
  assign T1795 = T1796 ^ 1'h1;
  assign T1796 = T1231 | T1239;
  assign readyToXmit_4_4 = T1797;
  assign T1797 = T1811 ? T1807 : T1798;
  assign T1798 = T1803 ? T1799 : 1'h0;
  assign T1799 = T1800 & RouterBuffer_4_io_deq_valid;
  assign T1800 = T1801 & T1021;
  assign T1801 = T1085 & T1802;
  assign T1802 = 3'h3 <= VCRouterStateManagement_4_io_currentState;
  assign T1803 = T1094 & T1804;
  assign T1804 = T1805[3'h4:3'h4];
  assign T1805 = 1'h1 << T1806;
  assign T1806 = R1015;
  assign T1807 = T1808 & RouterBuffer_4_io_deq_valid;
  assign T1808 = T1809 & T1021;
  assign T1809 = T1085 & T1810;
  assign T1810 = VCRouterStateManagement_4_io_currentState == 3'h4;
  assign T1811 = T1812 & T1804;
  assign T1812 = T1813 ^ 1'h1;
  assign T1813 = T1087 | T1095;
  assign T1814 = {T1868, T1815};
  assign T1815 = {readyToXmit_7_4, T1816};
  assign T1816 = {readyToXmit_6_4, readyToXmit_5_4};
  assign readyToXmit_5_4 = T1817;
  assign T1817 = T1831 ? T1827 : T1818;
  assign T1818 = T1823 ? T1819 : 1'h0;
  assign T1819 = T1820 & RouterBuffer_5_io_deq_valid;
  assign T1820 = T1821 & T877;
  assign T1821 = T941 & T1822;
  assign T1822 = 3'h3 <= VCRouterStateManagement_5_io_currentState;
  assign T1823 = T950 & T1824;
  assign T1824 = T1825[3'h4:3'h4];
  assign T1825 = 1'h1 << T1826;
  assign T1826 = R871;
  assign T1827 = T1828 & RouterBuffer_5_io_deq_valid;
  assign T1828 = T1829 & T877;
  assign T1829 = T941 & T1830;
  assign T1830 = VCRouterStateManagement_5_io_currentState == 3'h4;
  assign T1831 = T1832 & T1824;
  assign T1832 = T1833 ^ 1'h1;
  assign T1833 = T943 | T951;
  assign readyToXmit_6_4 = T1834;
  assign T1834 = T1848 ? T1844 : T1835;
  assign T1835 = T1840 ? T1836 : 1'h0;
  assign T1836 = T1837 & RouterBuffer_6_io_deq_valid;
  assign T1837 = T1838 & T733;
  assign T1838 = T797 & T1839;
  assign T1839 = 3'h3 <= VCRouterStateManagement_6_io_currentState;
  assign T1840 = T806 & T1841;
  assign T1841 = T1842[3'h4:3'h4];
  assign T1842 = 1'h1 << T1843;
  assign T1843 = R727;
  assign T1844 = T1845 & RouterBuffer_6_io_deq_valid;
  assign T1845 = T1846 & T733;
  assign T1846 = T797 & T1847;
  assign T1847 = VCRouterStateManagement_6_io_currentState == 3'h4;
  assign T1848 = T1849 & T1841;
  assign T1849 = T1850 ^ 1'h1;
  assign T1850 = T799 | T807;
  assign readyToXmit_7_4 = T1851;
  assign T1851 = T1865 ? T1861 : T1852;
  assign T1852 = T1857 ? T1853 : 1'h0;
  assign T1853 = T1854 & RouterBuffer_7_io_deq_valid;
  assign T1854 = T1855 & T589;
  assign T1855 = T653 & T1856;
  assign T1856 = 3'h3 <= VCRouterStateManagement_7_io_currentState;
  assign T1857 = T662 & T1858;
  assign T1858 = T1859[3'h4:3'h4];
  assign T1859 = 1'h1 << T1860;
  assign T1860 = R583;
  assign T1861 = T1862 & RouterBuffer_7_io_deq_valid;
  assign T1862 = T1863 & T589;
  assign T1863 = T653 & T1864;
  assign T1864 = VCRouterStateManagement_7_io_currentState == 3'h4;
  assign T1865 = T1866 & T1858;
  assign T1866 = T1867 ^ 1'h1;
  assign T1867 = T655 | T663;
  assign T1868 = {readyToXmit_9_4, readyToXmit_8_4};
  assign readyToXmit_8_4 = T1869;
  assign T1869 = T1883 ? T1879 : T1870;
  assign T1870 = T1875 ? T1871 : 1'h0;
  assign T1871 = T1872 & RouterBuffer_8_io_deq_valid;
  assign T1872 = T1873 & T445;
  assign T1873 = T509 & T1874;
  assign T1874 = 3'h3 <= VCRouterStateManagement_8_io_currentState;
  assign T1875 = T518 & T1876;
  assign T1876 = T1877[3'h4:3'h4];
  assign T1877 = 1'h1 << T1878;
  assign T1878 = R439;
  assign T1879 = T1880 & RouterBuffer_8_io_deq_valid;
  assign T1880 = T1881 & T445;
  assign T1881 = T509 & T1882;
  assign T1882 = VCRouterStateManagement_8_io_currentState == 3'h4;
  assign T1883 = T1884 & T1876;
  assign T1884 = T1885 ^ 1'h1;
  assign T1885 = T511 | T519;
  assign readyToXmit_9_4 = T1886;
  assign T1886 = T1900 ? T1896 : T1887;
  assign T1887 = T1892 ? T1888 : 1'h0;
  assign T1888 = T1889 & RouterBuffer_9_io_deq_valid;
  assign T1889 = T1890 & T301;
  assign T1890 = T365 & T1891;
  assign T1891 = 3'h3 <= VCRouterStateManagement_9_io_currentState;
  assign T1892 = T374 & T1893;
  assign T1893 = T1894[3'h4:3'h4];
  assign T1894 = 1'h1 << T1895;
  assign T1895 = R295;
  assign T1896 = T1897 & RouterBuffer_9_io_deq_valid;
  assign T1897 = T1898 & T301;
  assign T1898 = T365 & T1899;
  assign T1899 = VCRouterStateManagement_9_io_currentState == 3'h4;
  assign T1900 = T1901 & T1893;
  assign T1901 = T1902 ^ 1'h1;
  assign T1902 = T367 | T375;
  assign T1903 = T1904 ? CreditCon_7_io_outCredit : CreditCon_6_io_outCredit;
  assign T1904 = T234;
  assign T1905 = T1906 != 10'h0;
  assign T1906 = T1907;
  assign T1907 = {T1937, T1908};
  assign T1908 = {T1926, T1909};
  assign T1909 = {readyToXmit_2_3, T1910};
  assign T1910 = {readyToXmit_1_3, readyToXmit_0_3};
  assign readyToXmit_0_3 = T1911;
  assign T1911 = T1915 ? T1738 : T1912;
  assign T1912 = T1913 ? T1730 : 1'h0;
  assign T1913 = T1670 & T1914;
  assign T1914 = T1736[2'h3:2'h3];
  assign T1915 = T1743 & T1914;
  assign readyToXmit_1_3 = T1916;
  assign T1916 = T1920 ? T1755 : T1917;
  assign T1917 = T1918 ? T1747 : 1'h0;
  assign T1918 = T1526 & T1919;
  assign T1919 = T1753[2'h3:2'h3];
  assign T1920 = T1760 & T1919;
  assign readyToXmit_2_3 = T1921;
  assign T1921 = T1925 ? T1772 : T1922;
  assign T1922 = T1923 ? T1764 : 1'h0;
  assign T1923 = T1382 & T1924;
  assign T1924 = T1770[2'h3:2'h3];
  assign T1925 = T1777 & T1924;
  assign T1926 = {readyToXmit_4_3, readyToXmit_3_3};
  assign readyToXmit_3_3 = T1927;
  assign T1927 = T1931 ? T1790 : T1928;
  assign T1928 = T1929 ? T1782 : 1'h0;
  assign T1929 = T1238 & T1930;
  assign T1930 = T1788[2'h3:2'h3];
  assign T1931 = T1795 & T1930;
  assign readyToXmit_4_3 = T1932;
  assign T1932 = T1936 ? T1807 : T1933;
  assign T1933 = T1934 ? T1799 : 1'h0;
  assign T1934 = T1094 & T1935;
  assign T1935 = T1805[2'h3:2'h3];
  assign T1936 = T1812 & T1935;
  assign T1937 = {T1955, T1938};
  assign T1938 = {readyToXmit_7_3, T1939};
  assign T1939 = {readyToXmit_6_3, readyToXmit_5_3};
  assign readyToXmit_5_3 = T1940;
  assign T1940 = T1944 ? T1827 : T1941;
  assign T1941 = T1942 ? T1819 : 1'h0;
  assign T1942 = T950 & T1943;
  assign T1943 = T1825[2'h3:2'h3];
  assign T1944 = T1832 & T1943;
  assign readyToXmit_6_3 = T1945;
  assign T1945 = T1949 ? T1844 : T1946;
  assign T1946 = T1947 ? T1836 : 1'h0;
  assign T1947 = T806 & T1948;
  assign T1948 = T1842[2'h3:2'h3];
  assign T1949 = T1849 & T1948;
  assign readyToXmit_7_3 = T1950;
  assign T1950 = T1954 ? T1861 : T1951;
  assign T1951 = T1952 ? T1853 : 1'h0;
  assign T1952 = T662 & T1953;
  assign T1953 = T1859[2'h3:2'h3];
  assign T1954 = T1866 & T1953;
  assign T1955 = {readyToXmit_9_3, readyToXmit_8_3};
  assign readyToXmit_8_3 = T1956;
  assign T1956 = T1960 ? T1879 : T1957;
  assign T1957 = T1958 ? T1871 : 1'h0;
  assign T1958 = T518 & T1959;
  assign T1959 = T1877[2'h3:2'h3];
  assign T1960 = T1884 & T1959;
  assign readyToXmit_9_3 = T1961;
  assign T1961 = T1965 ? T1896 : T1962;
  assign T1962 = T1963 ? T1888 : 1'h0;
  assign T1963 = T374 & T1964;
  assign T1964 = T1894[2'h3:2'h3];
  assign T1965 = T1901 & T1964;
  assign T1966 = T1967 ? CreditCon_5_io_outCredit : CreditCon_4_io_outCredit;
  assign T1967 = T246;
  assign T1968 = T1969 != 10'h0;
  assign T1969 = T1970;
  assign T1970 = {T2000, T1971};
  assign T1971 = {T1989, T1972};
  assign T1972 = {readyToXmit_2_2, T1973};
  assign T1973 = {readyToXmit_1_2, readyToXmit_0_2};
  assign readyToXmit_0_2 = T1974;
  assign T1974 = T1978 ? T1738 : T1975;
  assign T1975 = T1976 ? T1730 : 1'h0;
  assign T1976 = T1670 & T1977;
  assign T1977 = T1736[2'h2:2'h2];
  assign T1978 = T1743 & T1977;
  assign readyToXmit_1_2 = T1979;
  assign T1979 = T1983 ? T1755 : T1980;
  assign T1980 = T1981 ? T1747 : 1'h0;
  assign T1981 = T1526 & T1982;
  assign T1982 = T1753[2'h2:2'h2];
  assign T1983 = T1760 & T1982;
  assign readyToXmit_2_2 = T1984;
  assign T1984 = T1988 ? T1772 : T1985;
  assign T1985 = T1986 ? T1764 : 1'h0;
  assign T1986 = T1382 & T1987;
  assign T1987 = T1770[2'h2:2'h2];
  assign T1988 = T1777 & T1987;
  assign T1989 = {readyToXmit_4_2, readyToXmit_3_2};
  assign readyToXmit_3_2 = T1990;
  assign T1990 = T1994 ? T1790 : T1991;
  assign T1991 = T1992 ? T1782 : 1'h0;
  assign T1992 = T1238 & T1993;
  assign T1993 = T1788[2'h2:2'h2];
  assign T1994 = T1795 & T1993;
  assign readyToXmit_4_2 = T1995;
  assign T1995 = T1999 ? T1807 : T1996;
  assign T1996 = T1997 ? T1799 : 1'h0;
  assign T1997 = T1094 & T1998;
  assign T1998 = T1805[2'h2:2'h2];
  assign T1999 = T1812 & T1998;
  assign T2000 = {T2018, T2001};
  assign T2001 = {readyToXmit_7_2, T2002};
  assign T2002 = {readyToXmit_6_2, readyToXmit_5_2};
  assign readyToXmit_5_2 = T2003;
  assign T2003 = T2007 ? T1827 : T2004;
  assign T2004 = T2005 ? T1819 : 1'h0;
  assign T2005 = T950 & T2006;
  assign T2006 = T1825[2'h2:2'h2];
  assign T2007 = T1832 & T2006;
  assign readyToXmit_6_2 = T2008;
  assign T2008 = T2012 ? T1844 : T2009;
  assign T2009 = T2010 ? T1836 : 1'h0;
  assign T2010 = T806 & T2011;
  assign T2011 = T1842[2'h2:2'h2];
  assign T2012 = T1849 & T2011;
  assign readyToXmit_7_2 = T2013;
  assign T2013 = T2017 ? T1861 : T2014;
  assign T2014 = T2015 ? T1853 : 1'h0;
  assign T2015 = T662 & T2016;
  assign T2016 = T1859[2'h2:2'h2];
  assign T2017 = T1866 & T2016;
  assign T2018 = {readyToXmit_9_2, readyToXmit_8_2};
  assign readyToXmit_8_2 = T2019;
  assign T2019 = T2023 ? T1879 : T2020;
  assign T2020 = T2021 ? T1871 : 1'h0;
  assign T2021 = T518 & T2022;
  assign T2022 = T1877[2'h2:2'h2];
  assign T2023 = T1884 & T2022;
  assign readyToXmit_9_2 = T2024;
  assign T2024 = T2028 ? T1896 : T2025;
  assign T2025 = T2026 ? T1888 : 1'h0;
  assign T2026 = T374 & T2027;
  assign T2027 = T1894[2'h2:2'h2];
  assign T2028 = T1901 & T2027;
  assign T2029 = T2030 ? CreditCon_3_io_outCredit : CreditCon_2_io_outCredit;
  assign T2030 = T258;
  assign T2031 = T2032 != 10'h0;
  assign T2032 = T2033;
  assign T2033 = {T2063, T2034};
  assign T2034 = {T2052, T2035};
  assign T2035 = {readyToXmit_2_1, T2036};
  assign T2036 = {readyToXmit_1_1, readyToXmit_0_1};
  assign readyToXmit_0_1 = T2037;
  assign T2037 = T2041 ? T1738 : T2038;
  assign T2038 = T2039 ? T1730 : 1'h0;
  assign T2039 = T1670 & T2040;
  assign T2040 = T1736[1'h1:1'h1];
  assign T2041 = T1743 & T2040;
  assign readyToXmit_1_1 = T2042;
  assign T2042 = T2046 ? T1755 : T2043;
  assign T2043 = T2044 ? T1747 : 1'h0;
  assign T2044 = T1526 & T2045;
  assign T2045 = T1753[1'h1:1'h1];
  assign T2046 = T1760 & T2045;
  assign readyToXmit_2_1 = T2047;
  assign T2047 = T2051 ? T1772 : T2048;
  assign T2048 = T2049 ? T1764 : 1'h0;
  assign T2049 = T1382 & T2050;
  assign T2050 = T1770[1'h1:1'h1];
  assign T2051 = T1777 & T2050;
  assign T2052 = {readyToXmit_4_1, readyToXmit_3_1};
  assign readyToXmit_3_1 = T2053;
  assign T2053 = T2057 ? T1790 : T2054;
  assign T2054 = T2055 ? T1782 : 1'h0;
  assign T2055 = T1238 & T2056;
  assign T2056 = T1788[1'h1:1'h1];
  assign T2057 = T1795 & T2056;
  assign readyToXmit_4_1 = T2058;
  assign T2058 = T2062 ? T1807 : T2059;
  assign T2059 = T2060 ? T1799 : 1'h0;
  assign T2060 = T1094 & T2061;
  assign T2061 = T1805[1'h1:1'h1];
  assign T2062 = T1812 & T2061;
  assign T2063 = {T2081, T2064};
  assign T2064 = {readyToXmit_7_1, T2065};
  assign T2065 = {readyToXmit_6_1, readyToXmit_5_1};
  assign readyToXmit_5_1 = T2066;
  assign T2066 = T2070 ? T1827 : T2067;
  assign T2067 = T2068 ? T1819 : 1'h0;
  assign T2068 = T950 & T2069;
  assign T2069 = T1825[1'h1:1'h1];
  assign T2070 = T1832 & T2069;
  assign readyToXmit_6_1 = T2071;
  assign T2071 = T2075 ? T1844 : T2072;
  assign T2072 = T2073 ? T1836 : 1'h0;
  assign T2073 = T806 & T2074;
  assign T2074 = T1842[1'h1:1'h1];
  assign T2075 = T1849 & T2074;
  assign readyToXmit_7_1 = T2076;
  assign T2076 = T2080 ? T1861 : T2077;
  assign T2077 = T2078 ? T1853 : 1'h0;
  assign T2078 = T662 & T2079;
  assign T2079 = T1859[1'h1:1'h1];
  assign T2080 = T1866 & T2079;
  assign T2081 = {readyToXmit_9_1, readyToXmit_8_1};
  assign readyToXmit_8_1 = T2082;
  assign T2082 = T2086 ? T1879 : T2083;
  assign T2083 = T2084 ? T1871 : 1'h0;
  assign T2084 = T518 & T2085;
  assign T2085 = T1877[1'h1:1'h1];
  assign T2086 = T1884 & T2085;
  assign readyToXmit_9_1 = T2087;
  assign T2087 = T2091 ? T1896 : T2088;
  assign T2088 = T2089 ? T1888 : 1'h0;
  assign T2089 = T374 & T2090;
  assign T2090 = T1894[1'h1:1'h1];
  assign T2091 = T1901 & T2090;
  assign T2092 = T2093 ? CreditCon_1_io_outCredit : CreditCon_io_outCredit;
  assign T2093 = T270;
  assign T2094 = T2095 != 10'h0;
  assign T2095 = T2096;
  assign T2096 = {T2126, T2097};
  assign T2097 = {T2115, T2098};
  assign T2098 = {readyToXmit_2_0, T2099};
  assign T2099 = {readyToXmit_1_0, readyToXmit_0_0};
  assign readyToXmit_0_0 = T2100;
  assign T2100 = T2104 ? T1738 : T2101;
  assign T2101 = T2102 ? T1730 : 1'h0;
  assign T2102 = T1670 & T2103;
  assign T2103 = T1736[1'h0:1'h0];
  assign T2104 = T1743 & T2103;
  assign readyToXmit_1_0 = T2105;
  assign T2105 = T2109 ? T1755 : T2106;
  assign T2106 = T2107 ? T1747 : 1'h0;
  assign T2107 = T1526 & T2108;
  assign T2108 = T1753[1'h0:1'h0];
  assign T2109 = T1760 & T2108;
  assign readyToXmit_2_0 = T2110;
  assign T2110 = T2114 ? T1772 : T2111;
  assign T2111 = T2112 ? T1764 : 1'h0;
  assign T2112 = T1382 & T2113;
  assign T2113 = T1770[1'h0:1'h0];
  assign T2114 = T1777 & T2113;
  assign T2115 = {readyToXmit_4_0, readyToXmit_3_0};
  assign readyToXmit_3_0 = T2116;
  assign T2116 = T2120 ? T1790 : T2117;
  assign T2117 = T2118 ? T1782 : 1'h0;
  assign T2118 = T1238 & T2119;
  assign T2119 = T1788[1'h0:1'h0];
  assign T2120 = T1795 & T2119;
  assign readyToXmit_4_0 = T2121;
  assign T2121 = T2125 ? T1807 : T2122;
  assign T2122 = T2123 ? T1799 : 1'h0;
  assign T2123 = T1094 & T2124;
  assign T2124 = T1805[1'h0:1'h0];
  assign T2125 = T1812 & T2124;
  assign T2126 = {T2144, T2127};
  assign T2127 = {readyToXmit_7_0, T2128};
  assign T2128 = {readyToXmit_6_0, readyToXmit_5_0};
  assign readyToXmit_5_0 = T2129;
  assign T2129 = T2133 ? T1827 : T2130;
  assign T2130 = T2131 ? T1819 : 1'h0;
  assign T2131 = T950 & T2132;
  assign T2132 = T1825[1'h0:1'h0];
  assign T2133 = T1832 & T2132;
  assign readyToXmit_6_0 = T2134;
  assign T2134 = T2138 ? T1844 : T2135;
  assign T2135 = T2136 ? T1836 : 1'h0;
  assign T2136 = T806 & T2137;
  assign T2137 = T1842[1'h0:1'h0];
  assign T2138 = T1849 & T2137;
  assign readyToXmit_7_0 = T2139;
  assign T2139 = T2143 ? T1861 : T2140;
  assign T2140 = T2141 ? T1853 : 1'h0;
  assign T2141 = T662 & T2142;
  assign T2142 = T1859[1'h0:1'h0];
  assign T2143 = T1866 & T2142;
  assign T2144 = {readyToXmit_9_0, readyToXmit_8_0};
  assign readyToXmit_8_0 = T2145;
  assign T2145 = T2149 ? T1879 : T2146;
  assign T2146 = T2147 ? T1871 : 1'h0;
  assign T2147 = T518 & T2148;
  assign T2148 = T1877[1'h0:1'h0];
  assign T2149 = T1884 & T2148;
  assign readyToXmit_9_0 = T2150;
  assign T2150 = T2154 ? T1896 : T2151;
  assign T2151 = T2152 ? T1888 : 1'h0;
  assign T2152 = T374 & T2153;
  assign T2153 = T1894[1'h0:1'h0];
  assign T2154 = T1901 & T2153;
  assign T2155 = RouterBuffer_io_deq_valid & T2156;
  assign T2156 = 3'h2 <= VCRouterStateManagement_io_currentState;
  assign T2157 = RouterBuffer_1_io_deq_valid & T2158;
  assign T2158 = 3'h2 <= VCRouterStateManagement_1_io_currentState;
  assign T2159 = RouterBuffer_2_io_deq_valid & T2160;
  assign T2160 = 3'h2 <= VCRouterStateManagement_2_io_currentState;
  assign T2161 = RouterBuffer_3_io_deq_valid & T2162;
  assign T2162 = 3'h2 <= VCRouterStateManagement_3_io_currentState;
  assign T2163 = RouterBuffer_4_io_deq_valid & T2164;
  assign T2164 = 3'h2 <= VCRouterStateManagement_4_io_currentState;
  assign T2165 = RouterBuffer_5_io_deq_valid & T2166;
  assign T2166 = 3'h2 <= VCRouterStateManagement_5_io_currentState;
  assign T2167 = RouterBuffer_6_io_deq_valid & T2168;
  assign T2168 = 3'h2 <= VCRouterStateManagement_6_io_currentState;
  assign T2169 = RouterBuffer_7_io_deq_valid & T2170;
  assign T2170 = 3'h2 <= VCRouterStateManagement_7_io_currentState;
  assign T2171 = RouterBuffer_8_io_deq_valid & T2172;
  assign T2172 = 3'h2 <= VCRouterStateManagement_8_io_currentState;
  assign T2173 = RouterBuffer_9_io_deq_valid & T2174;
  assign T2174 = 3'h2 <= VCRouterStateManagement_9_io_currentState;
  assign T2175 = validVCs_0_0[1'h0:1'h0];
  assign T2177 = T2179 & T2178;
  assign T2178 = VCRouterOutputStateManagement_io_currentState == 2'h2;
  assign T2179 = flitsAreTail_0 & CreditCon_io_outCredit;
  assign T2180 = validVCs_0_0[1'h1:1'h1];
  assign T2182 = T2184 & T2183;
  assign T2183 = VCRouterOutputStateManagement_io_currentState == 2'h2;
  assign T2184 = flitsAreTail_0 & CreditCon_1_io_outCredit;
  assign T2185 = validVCs_0_1[1'h0:1'h0];
  assign T2187 = T2189 & T2188;
  assign T2188 = VCRouterOutputStateManagement_1_io_currentState == 2'h2;
  assign T2189 = flitsAreTail_0 & CreditCon_2_io_outCredit;
  assign T2190 = validVCs_0_1[1'h1:1'h1];
  assign T2192 = T2194 & T2193;
  assign T2193 = VCRouterOutputStateManagement_1_io_currentState == 2'h2;
  assign T2194 = flitsAreTail_0 & CreditCon_3_io_outCredit;
  assign T2195 = validVCs_0_2[1'h0:1'h0];
  assign T2197 = T2199 & T2198;
  assign T2198 = VCRouterOutputStateManagement_2_io_currentState == 2'h2;
  assign T2199 = flitsAreTail_0 & CreditCon_4_io_outCredit;
  assign T2200 = validVCs_0_2[1'h1:1'h1];
  assign T2202 = T2204 & T2203;
  assign T2203 = VCRouterOutputStateManagement_2_io_currentState == 2'h2;
  assign T2204 = flitsAreTail_0 & CreditCon_5_io_outCredit;
  assign T2205 = validVCs_0_3[1'h0:1'h0];
  assign T2207 = T2209 & T2208;
  assign T2208 = VCRouterOutputStateManagement_3_io_currentState == 2'h2;
  assign T2209 = flitsAreTail_0 & CreditCon_6_io_outCredit;
  assign T2210 = validVCs_0_3[1'h1:1'h1];
  assign T2212 = T2214 & T2213;
  assign T2213 = VCRouterOutputStateManagement_3_io_currentState == 2'h2;
  assign T2214 = flitsAreTail_0 & CreditCon_7_io_outCredit;
  assign T2215 = validVCs_0_4[1'h0:1'h0];
  assign T2217 = T2219 & T2218;
  assign T2218 = VCRouterOutputStateManagement_4_io_currentState == 2'h2;
  assign T2219 = flitsAreTail_0 & CreditCon_8_io_outCredit;
  assign T2220 = validVCs_0_4[1'h1:1'h1];
  assign T2222 = T2224 & T2223;
  assign T2223 = VCRouterOutputStateManagement_4_io_currentState == 2'h2;
  assign T2224 = flitsAreTail_0 & CreditCon_9_io_outCredit;
  assign T2225 = validVCs_1_0[1'h0:1'h0];
  assign T2227 = T2229 & T2228;
  assign T2228 = VCRouterOutputStateManagement_io_currentState == 2'h2;
  assign T2229 = flitsAreTail_1 & CreditCon_io_outCredit;
  assign T2230 = validVCs_1_0[1'h1:1'h1];
  assign T2232 = T2234 & T2233;
  assign T2233 = VCRouterOutputStateManagement_io_currentState == 2'h2;
  assign T2234 = flitsAreTail_1 & CreditCon_1_io_outCredit;
  assign T2235 = validVCs_1_1[1'h0:1'h0];
  assign T2237 = T2239 & T2238;
  assign T2238 = VCRouterOutputStateManagement_1_io_currentState == 2'h2;
  assign T2239 = flitsAreTail_1 & CreditCon_2_io_outCredit;
  assign T2240 = validVCs_1_1[1'h1:1'h1];
  assign T2242 = T2244 & T2243;
  assign T2243 = VCRouterOutputStateManagement_1_io_currentState == 2'h2;
  assign T2244 = flitsAreTail_1 & CreditCon_3_io_outCredit;
  assign T2245 = validVCs_1_2[1'h0:1'h0];
  assign T2247 = T2249 & T2248;
  assign T2248 = VCRouterOutputStateManagement_2_io_currentState == 2'h2;
  assign T2249 = flitsAreTail_1 & CreditCon_4_io_outCredit;
  assign T2250 = validVCs_1_2[1'h1:1'h1];
  assign T2252 = T2254 & T2253;
  assign T2253 = VCRouterOutputStateManagement_2_io_currentState == 2'h2;
  assign T2254 = flitsAreTail_1 & CreditCon_5_io_outCredit;
  assign T2255 = validVCs_1_3[1'h0:1'h0];
  assign T2257 = T2259 & T2258;
  assign T2258 = VCRouterOutputStateManagement_3_io_currentState == 2'h2;
  assign T2259 = flitsAreTail_1 & CreditCon_6_io_outCredit;
  assign T2260 = validVCs_1_3[1'h1:1'h1];
  assign T2262 = T2264 & T2263;
  assign T2263 = VCRouterOutputStateManagement_3_io_currentState == 2'h2;
  assign T2264 = flitsAreTail_1 & CreditCon_7_io_outCredit;
  assign T2265 = validVCs_1_4[1'h0:1'h0];
  assign T2267 = T2269 & T2268;
  assign T2268 = VCRouterOutputStateManagement_4_io_currentState == 2'h2;
  assign T2269 = flitsAreTail_1 & CreditCon_8_io_outCredit;
  assign T2270 = validVCs_1_4[1'h1:1'h1];
  assign T2272 = T2274 & T2273;
  assign T2273 = VCRouterOutputStateManagement_4_io_currentState == 2'h2;
  assign T2274 = flitsAreTail_1 & CreditCon_9_io_outCredit;
  assign T2275 = validVCs_2_0[1'h0:1'h0];
  assign T2277 = T2279 & T2278;
  assign T2278 = VCRouterOutputStateManagement_io_currentState == 2'h2;
  assign T2279 = flitsAreTail_2 & CreditCon_io_outCredit;
  assign T2280 = validVCs_2_0[1'h1:1'h1];
  assign T2282 = T2284 & T2283;
  assign T2283 = VCRouterOutputStateManagement_io_currentState == 2'h2;
  assign T2284 = flitsAreTail_2 & CreditCon_1_io_outCredit;
  assign T2285 = validVCs_2_1[1'h0:1'h0];
  assign T2287 = T2289 & T2288;
  assign T2288 = VCRouterOutputStateManagement_1_io_currentState == 2'h2;
  assign T2289 = flitsAreTail_2 & CreditCon_2_io_outCredit;
  assign T2290 = validVCs_2_1[1'h1:1'h1];
  assign T2292 = T2294 & T2293;
  assign T2293 = VCRouterOutputStateManagement_1_io_currentState == 2'h2;
  assign T2294 = flitsAreTail_2 & CreditCon_3_io_outCredit;
  assign T2295 = validVCs_2_2[1'h0:1'h0];
  assign T2297 = T2299 & T2298;
  assign T2298 = VCRouterOutputStateManagement_2_io_currentState == 2'h2;
  assign T2299 = flitsAreTail_2 & CreditCon_4_io_outCredit;
  assign T2300 = validVCs_2_2[1'h1:1'h1];
  assign T2302 = T2304 & T2303;
  assign T2303 = VCRouterOutputStateManagement_2_io_currentState == 2'h2;
  assign T2304 = flitsAreTail_2 & CreditCon_5_io_outCredit;
  assign T2305 = validVCs_2_3[1'h0:1'h0];
  assign T2307 = T2309 & T2308;
  assign T2308 = VCRouterOutputStateManagement_3_io_currentState == 2'h2;
  assign T2309 = flitsAreTail_2 & CreditCon_6_io_outCredit;
  assign T2310 = validVCs_2_3[1'h1:1'h1];
  assign T2312 = T2314 & T2313;
  assign T2313 = VCRouterOutputStateManagement_3_io_currentState == 2'h2;
  assign T2314 = flitsAreTail_2 & CreditCon_7_io_outCredit;
  assign T2315 = validVCs_2_4[1'h0:1'h0];
  assign T2317 = T2319 & T2318;
  assign T2318 = VCRouterOutputStateManagement_4_io_currentState == 2'h2;
  assign T2319 = flitsAreTail_2 & CreditCon_8_io_outCredit;
  assign T2320 = validVCs_2_4[1'h1:1'h1];
  assign T2322 = T2324 & T2323;
  assign T2323 = VCRouterOutputStateManagement_4_io_currentState == 2'h2;
  assign T2324 = flitsAreTail_2 & CreditCon_9_io_outCredit;
  assign T2325 = validVCs_3_0[1'h0:1'h0];
  assign T2327 = T2329 & T2328;
  assign T2328 = VCRouterOutputStateManagement_io_currentState == 2'h2;
  assign T2329 = flitsAreTail_3 & CreditCon_io_outCredit;
  assign T2330 = validVCs_3_0[1'h1:1'h1];
  assign T2332 = T2334 & T2333;
  assign T2333 = VCRouterOutputStateManagement_io_currentState == 2'h2;
  assign T2334 = flitsAreTail_3 & CreditCon_1_io_outCredit;
  assign T2335 = validVCs_3_1[1'h0:1'h0];
  assign T2337 = T2339 & T2338;
  assign T2338 = VCRouterOutputStateManagement_1_io_currentState == 2'h2;
  assign T2339 = flitsAreTail_3 & CreditCon_2_io_outCredit;
  assign T2340 = validVCs_3_1[1'h1:1'h1];
  assign T2342 = T2344 & T2343;
  assign T2343 = VCRouterOutputStateManagement_1_io_currentState == 2'h2;
  assign T2344 = flitsAreTail_3 & CreditCon_3_io_outCredit;
  assign T2345 = validVCs_3_2[1'h0:1'h0];
  assign T2347 = T2349 & T2348;
  assign T2348 = VCRouterOutputStateManagement_2_io_currentState == 2'h2;
  assign T2349 = flitsAreTail_3 & CreditCon_4_io_outCredit;
  assign T2350 = validVCs_3_2[1'h1:1'h1];
  assign T2352 = T2354 & T2353;
  assign T2353 = VCRouterOutputStateManagement_2_io_currentState == 2'h2;
  assign T2354 = flitsAreTail_3 & CreditCon_5_io_outCredit;
  assign T2355 = validVCs_3_3[1'h0:1'h0];
  assign T2357 = T2359 & T2358;
  assign T2358 = VCRouterOutputStateManagement_3_io_currentState == 2'h2;
  assign T2359 = flitsAreTail_3 & CreditCon_6_io_outCredit;
  assign T2360 = validVCs_3_3[1'h1:1'h1];
  assign T2362 = T2364 & T2363;
  assign T2363 = VCRouterOutputStateManagement_3_io_currentState == 2'h2;
  assign T2364 = flitsAreTail_3 & CreditCon_7_io_outCredit;
  assign T2365 = validVCs_3_4[1'h0:1'h0];
  assign T2367 = T2369 & T2368;
  assign T2368 = VCRouterOutputStateManagement_4_io_currentState == 2'h2;
  assign T2369 = flitsAreTail_3 & CreditCon_8_io_outCredit;
  assign T2370 = validVCs_3_4[1'h1:1'h1];
  assign T2372 = T2374 & T2373;
  assign T2373 = VCRouterOutputStateManagement_4_io_currentState == 2'h2;
  assign T2374 = flitsAreTail_3 & CreditCon_9_io_outCredit;
  assign T2375 = validVCs_4_0[1'h0:1'h0];
  assign T2377 = T2379 & T2378;
  assign T2378 = VCRouterOutputStateManagement_io_currentState == 2'h2;
  assign T2379 = flitsAreTail_4 & CreditCon_io_outCredit;
  assign T2380 = validVCs_4_0[1'h1:1'h1];
  assign T2382 = T2384 & T2383;
  assign T2383 = VCRouterOutputStateManagement_io_currentState == 2'h2;
  assign T2384 = flitsAreTail_4 & CreditCon_1_io_outCredit;
  assign T2385 = validVCs_4_1[1'h0:1'h0];
  assign T2387 = T2389 & T2388;
  assign T2388 = VCRouterOutputStateManagement_1_io_currentState == 2'h2;
  assign T2389 = flitsAreTail_4 & CreditCon_2_io_outCredit;
  assign T2390 = validVCs_4_1[1'h1:1'h1];
  assign T2392 = T2394 & T2393;
  assign T2393 = VCRouterOutputStateManagement_1_io_currentState == 2'h2;
  assign T2394 = flitsAreTail_4 & CreditCon_3_io_outCredit;
  assign T2395 = validVCs_4_2[1'h0:1'h0];
  assign T2397 = T2399 & T2398;
  assign T2398 = VCRouterOutputStateManagement_2_io_currentState == 2'h2;
  assign T2399 = flitsAreTail_4 & CreditCon_4_io_outCredit;
  assign T2400 = validVCs_4_2[1'h1:1'h1];
  assign T2402 = T2404 & T2403;
  assign T2403 = VCRouterOutputStateManagement_2_io_currentState == 2'h2;
  assign T2404 = flitsAreTail_4 & CreditCon_5_io_outCredit;
  assign T2405 = validVCs_4_3[1'h0:1'h0];
  assign T2407 = T2409 & T2408;
  assign T2408 = VCRouterOutputStateManagement_3_io_currentState == 2'h2;
  assign T2409 = flitsAreTail_4 & CreditCon_6_io_outCredit;
  assign T2410 = validVCs_4_3[1'h1:1'h1];
  assign T2412 = T2414 & T2413;
  assign T2413 = VCRouterOutputStateManagement_3_io_currentState == 2'h2;
  assign T2414 = flitsAreTail_4 & CreditCon_7_io_outCredit;
  assign T2415 = validVCs_4_4[1'h0:1'h0];
  assign T2417 = T2419 & T2418;
  assign T2418 = VCRouterOutputStateManagement_4_io_currentState == 2'h2;
  assign T2419 = flitsAreTail_4 & CreditCon_8_io_outCredit;
  assign T2420 = validVCs_4_4[1'h1:1'h1];
  assign T2422 = T2424 & T2423;
  assign T2423 = VCRouterOutputStateManagement_4_io_currentState == 2'h2;
  assign T2424 = flitsAreTail_4 & CreditCon_9_io_outCredit;
  assign T2425 = validVCs_5_0[1'h0:1'h0];
  assign T2427 = T2429 & T2428;
  assign T2428 = VCRouterOutputStateManagement_io_currentState == 2'h2;
  assign T2429 = flitsAreTail_5 & CreditCon_io_outCredit;
  assign T2430 = validVCs_5_0[1'h1:1'h1];
  assign T2432 = T2434 & T2433;
  assign T2433 = VCRouterOutputStateManagement_io_currentState == 2'h2;
  assign T2434 = flitsAreTail_5 & CreditCon_1_io_outCredit;
  assign T2435 = validVCs_5_1[1'h0:1'h0];
  assign T2437 = T2439 & T2438;
  assign T2438 = VCRouterOutputStateManagement_1_io_currentState == 2'h2;
  assign T2439 = flitsAreTail_5 & CreditCon_2_io_outCredit;
  assign T2440 = validVCs_5_1[1'h1:1'h1];
  assign T2442 = T2444 & T2443;
  assign T2443 = VCRouterOutputStateManagement_1_io_currentState == 2'h2;
  assign T2444 = flitsAreTail_5 & CreditCon_3_io_outCredit;
  assign T2445 = validVCs_5_2[1'h0:1'h0];
  assign T2447 = T2449 & T2448;
  assign T2448 = VCRouterOutputStateManagement_2_io_currentState == 2'h2;
  assign T2449 = flitsAreTail_5 & CreditCon_4_io_outCredit;
  assign T2450 = validVCs_5_2[1'h1:1'h1];
  assign T2452 = T2454 & T2453;
  assign T2453 = VCRouterOutputStateManagement_2_io_currentState == 2'h2;
  assign T2454 = flitsAreTail_5 & CreditCon_5_io_outCredit;
  assign T2455 = validVCs_5_3[1'h0:1'h0];
  assign T2457 = T2459 & T2458;
  assign T2458 = VCRouterOutputStateManagement_3_io_currentState == 2'h2;
  assign T2459 = flitsAreTail_5 & CreditCon_6_io_outCredit;
  assign T2460 = validVCs_5_3[1'h1:1'h1];
  assign T2462 = T2464 & T2463;
  assign T2463 = VCRouterOutputStateManagement_3_io_currentState == 2'h2;
  assign T2464 = flitsAreTail_5 & CreditCon_7_io_outCredit;
  assign T2465 = validVCs_5_4[1'h0:1'h0];
  assign T2467 = T2469 & T2468;
  assign T2468 = VCRouterOutputStateManagement_4_io_currentState == 2'h2;
  assign T2469 = flitsAreTail_5 & CreditCon_8_io_outCredit;
  assign T2470 = validVCs_5_4[1'h1:1'h1];
  assign T2472 = T2474 & T2473;
  assign T2473 = VCRouterOutputStateManagement_4_io_currentState == 2'h2;
  assign T2474 = flitsAreTail_5 & CreditCon_9_io_outCredit;
  assign T2475 = validVCs_6_0[1'h0:1'h0];
  assign T2477 = T2479 & T2478;
  assign T2478 = VCRouterOutputStateManagement_io_currentState == 2'h2;
  assign T2479 = flitsAreTail_6 & CreditCon_io_outCredit;
  assign T2480 = validVCs_6_0[1'h1:1'h1];
  assign T2482 = T2484 & T2483;
  assign T2483 = VCRouterOutputStateManagement_io_currentState == 2'h2;
  assign T2484 = flitsAreTail_6 & CreditCon_1_io_outCredit;
  assign T2485 = validVCs_6_1[1'h0:1'h0];
  assign T2487 = T2489 & T2488;
  assign T2488 = VCRouterOutputStateManagement_1_io_currentState == 2'h2;
  assign T2489 = flitsAreTail_6 & CreditCon_2_io_outCredit;
  assign T2490 = validVCs_6_1[1'h1:1'h1];
  assign T2492 = T2494 & T2493;
  assign T2493 = VCRouterOutputStateManagement_1_io_currentState == 2'h2;
  assign T2494 = flitsAreTail_6 & CreditCon_3_io_outCredit;
  assign T2495 = validVCs_6_2[1'h0:1'h0];
  assign T2497 = T2499 & T2498;
  assign T2498 = VCRouterOutputStateManagement_2_io_currentState == 2'h2;
  assign T2499 = flitsAreTail_6 & CreditCon_4_io_outCredit;
  assign T2500 = validVCs_6_2[1'h1:1'h1];
  assign T2502 = T2504 & T2503;
  assign T2503 = VCRouterOutputStateManagement_2_io_currentState == 2'h2;
  assign T2504 = flitsAreTail_6 & CreditCon_5_io_outCredit;
  assign T2505 = validVCs_6_3[1'h0:1'h0];
  assign T2507 = T2509 & T2508;
  assign T2508 = VCRouterOutputStateManagement_3_io_currentState == 2'h2;
  assign T2509 = flitsAreTail_6 & CreditCon_6_io_outCredit;
  assign T2510 = validVCs_6_3[1'h1:1'h1];
  assign T2512 = T2514 & T2513;
  assign T2513 = VCRouterOutputStateManagement_3_io_currentState == 2'h2;
  assign T2514 = flitsAreTail_6 & CreditCon_7_io_outCredit;
  assign T2515 = validVCs_6_4[1'h0:1'h0];
  assign T2517 = T2519 & T2518;
  assign T2518 = VCRouterOutputStateManagement_4_io_currentState == 2'h2;
  assign T2519 = flitsAreTail_6 & CreditCon_8_io_outCredit;
  assign T2520 = validVCs_6_4[1'h1:1'h1];
  assign T2522 = T2524 & T2523;
  assign T2523 = VCRouterOutputStateManagement_4_io_currentState == 2'h2;
  assign T2524 = flitsAreTail_6 & CreditCon_9_io_outCredit;
  assign T2525 = validVCs_7_0[1'h0:1'h0];
  assign T2527 = T2529 & T2528;
  assign T2528 = VCRouterOutputStateManagement_io_currentState == 2'h2;
  assign T2529 = flitsAreTail_7 & CreditCon_io_outCredit;
  assign T2530 = validVCs_7_0[1'h1:1'h1];
  assign T2532 = T2534 & T2533;
  assign T2533 = VCRouterOutputStateManagement_io_currentState == 2'h2;
  assign T2534 = flitsAreTail_7 & CreditCon_1_io_outCredit;
  assign T2535 = validVCs_7_1[1'h0:1'h0];
  assign T2537 = T2539 & T2538;
  assign T2538 = VCRouterOutputStateManagement_1_io_currentState == 2'h2;
  assign T2539 = flitsAreTail_7 & CreditCon_2_io_outCredit;
  assign T2540 = validVCs_7_1[1'h1:1'h1];
  assign T2542 = T2544 & T2543;
  assign T2543 = VCRouterOutputStateManagement_1_io_currentState == 2'h2;
  assign T2544 = flitsAreTail_7 & CreditCon_3_io_outCredit;
  assign T2545 = validVCs_7_2[1'h0:1'h0];
  assign T2547 = T2549 & T2548;
  assign T2548 = VCRouterOutputStateManagement_2_io_currentState == 2'h2;
  assign T2549 = flitsAreTail_7 & CreditCon_4_io_outCredit;
  assign T2550 = validVCs_7_2[1'h1:1'h1];
  assign T2552 = T2554 & T2553;
  assign T2553 = VCRouterOutputStateManagement_2_io_currentState == 2'h2;
  assign T2554 = flitsAreTail_7 & CreditCon_5_io_outCredit;
  assign T2555 = validVCs_7_3[1'h0:1'h0];
  assign T2557 = T2559 & T2558;
  assign T2558 = VCRouterOutputStateManagement_3_io_currentState == 2'h2;
  assign T2559 = flitsAreTail_7 & CreditCon_6_io_outCredit;
  assign T2560 = validVCs_7_3[1'h1:1'h1];
  assign T2562 = T2564 & T2563;
  assign T2563 = VCRouterOutputStateManagement_3_io_currentState == 2'h2;
  assign T2564 = flitsAreTail_7 & CreditCon_7_io_outCredit;
  assign T2565 = validVCs_7_4[1'h0:1'h0];
  assign T2567 = T2569 & T2568;
  assign T2568 = VCRouterOutputStateManagement_4_io_currentState == 2'h2;
  assign T2569 = flitsAreTail_7 & CreditCon_8_io_outCredit;
  assign T2570 = validVCs_7_4[1'h1:1'h1];
  assign T2572 = T2574 & T2573;
  assign T2573 = VCRouterOutputStateManagement_4_io_currentState == 2'h2;
  assign T2574 = flitsAreTail_7 & CreditCon_9_io_outCredit;
  assign T2575 = validVCs_8_0[1'h0:1'h0];
  assign T2577 = T2579 & T2578;
  assign T2578 = VCRouterOutputStateManagement_io_currentState == 2'h2;
  assign T2579 = flitsAreTail_8 & CreditCon_io_outCredit;
  assign T2580 = validVCs_8_0[1'h1:1'h1];
  assign T2582 = T2584 & T2583;
  assign T2583 = VCRouterOutputStateManagement_io_currentState == 2'h2;
  assign T2584 = flitsAreTail_8 & CreditCon_1_io_outCredit;
  assign T2585 = validVCs_8_1[1'h0:1'h0];
  assign T2587 = T2589 & T2588;
  assign T2588 = VCRouterOutputStateManagement_1_io_currentState == 2'h2;
  assign T2589 = flitsAreTail_8 & CreditCon_2_io_outCredit;
  assign T2590 = validVCs_8_1[1'h1:1'h1];
  assign T2592 = T2594 & T2593;
  assign T2593 = VCRouterOutputStateManagement_1_io_currentState == 2'h2;
  assign T2594 = flitsAreTail_8 & CreditCon_3_io_outCredit;
  assign T2595 = validVCs_8_2[1'h0:1'h0];
  assign T2597 = T2599 & T2598;
  assign T2598 = VCRouterOutputStateManagement_2_io_currentState == 2'h2;
  assign T2599 = flitsAreTail_8 & CreditCon_4_io_outCredit;
  assign T2600 = validVCs_8_2[1'h1:1'h1];
  assign T2602 = T2604 & T2603;
  assign T2603 = VCRouterOutputStateManagement_2_io_currentState == 2'h2;
  assign T2604 = flitsAreTail_8 & CreditCon_5_io_outCredit;
  assign T2605 = validVCs_8_3[1'h0:1'h0];
  assign T2607 = T2609 & T2608;
  assign T2608 = VCRouterOutputStateManagement_3_io_currentState == 2'h2;
  assign T2609 = flitsAreTail_8 & CreditCon_6_io_outCredit;
  assign T2610 = validVCs_8_3[1'h1:1'h1];
  assign T2612 = T2614 & T2613;
  assign T2613 = VCRouterOutputStateManagement_3_io_currentState == 2'h2;
  assign T2614 = flitsAreTail_8 & CreditCon_7_io_outCredit;
  assign T2615 = validVCs_8_4[1'h0:1'h0];
  assign T2617 = T2619 & T2618;
  assign T2618 = VCRouterOutputStateManagement_4_io_currentState == 2'h2;
  assign T2619 = flitsAreTail_8 & CreditCon_8_io_outCredit;
  assign T2620 = validVCs_8_4[1'h1:1'h1];
  assign T2622 = T2624 & T2623;
  assign T2623 = VCRouterOutputStateManagement_4_io_currentState == 2'h2;
  assign T2624 = flitsAreTail_8 & CreditCon_9_io_outCredit;
  assign T2625 = validVCs_9_0[1'h0:1'h0];
  assign T2627 = T2629 & T2628;
  assign T2628 = VCRouterOutputStateManagement_io_currentState == 2'h2;
  assign T2629 = flitsAreTail_9 & CreditCon_io_outCredit;
  assign T2630 = validVCs_9_0[1'h1:1'h1];
  assign T2632 = T2634 & T2633;
  assign T2633 = VCRouterOutputStateManagement_io_currentState == 2'h2;
  assign T2634 = flitsAreTail_9 & CreditCon_1_io_outCredit;
  assign T2635 = validVCs_9_1[1'h0:1'h0];
  assign T2637 = T2639 & T2638;
  assign T2638 = VCRouterOutputStateManagement_1_io_currentState == 2'h2;
  assign T2639 = flitsAreTail_9 & CreditCon_2_io_outCredit;
  assign T2640 = validVCs_9_1[1'h1:1'h1];
  assign T2642 = T2644 & T2643;
  assign T2643 = VCRouterOutputStateManagement_1_io_currentState == 2'h2;
  assign T2644 = flitsAreTail_9 & CreditCon_3_io_outCredit;
  assign T2645 = validVCs_9_2[1'h0:1'h0];
  assign T2647 = T2649 & T2648;
  assign T2648 = VCRouterOutputStateManagement_2_io_currentState == 2'h2;
  assign T2649 = flitsAreTail_9 & CreditCon_4_io_outCredit;
  assign T2650 = validVCs_9_2[1'h1:1'h1];
  assign T2652 = T2654 & T2653;
  assign T2653 = VCRouterOutputStateManagement_2_io_currentState == 2'h2;
  assign T2654 = flitsAreTail_9 & CreditCon_5_io_outCredit;
  assign T2655 = validVCs_9_3[1'h0:1'h0];
  assign T2657 = T2659 & T2658;
  assign T2658 = VCRouterOutputStateManagement_3_io_currentState == 2'h2;
  assign T2659 = flitsAreTail_9 & CreditCon_6_io_outCredit;
  assign T2660 = validVCs_9_3[1'h1:1'h1];
  assign T2662 = T2664 & T2663;
  assign T2663 = VCRouterOutputStateManagement_3_io_currentState == 2'h2;
  assign T2664 = flitsAreTail_9 & CreditCon_7_io_outCredit;
  assign T2665 = validVCs_9_4[1'h0:1'h0];
  assign T2667 = T2669 & T2668;
  assign T2668 = VCRouterOutputStateManagement_4_io_currentState == 2'h2;
  assign T2669 = flitsAreTail_9 & CreditCon_8_io_outCredit;
  assign T2670 = validVCs_9_4[1'h1:1'h1];
  assign T2672 = T2674 & T2673;
  assign T2673 = VCRouterOutputStateManagement_4_io_currentState == 2'h2;
  assign T2674 = flitsAreTail_9 & CreditCon_9_io_outCredit;
  assign T3182 = reset ? 3'h0 : T2676;
  assign T2676 = T1670 ? T2677 : R2675;
  assign T2677 = T2678[2'h2:1'h0];
  assign T2678 = RouterBuffer_io_deq_bits_x[5'h1f:1'h1];
  assign T2679 = T2681 & T2680;
  assign T2680 = 3'h3 <= VCRouterStateManagement_io_currentState;
  assign T2681 = T2682;
  assign T2682 = R2683[1'h0:1'h0];
  assign T3183 = reset ? 8'h0 : T2684;
  assign T2684 = 1'h1 << CMeshDOR_io_result;
  assign T2685 = T2687 & T2686;
  assign T2686 = VCRouterStateManagement_io_currentState == 3'h4;
  assign T2687 = R2688;
  assign T3184 = reset ? 1'h1 : T1692;
  assign T3185 = reset ? 3'h0 : T2690;
  assign T2690 = T1526 ? T2691 : R2689;
  assign T2691 = T2692[2'h2:1'h0];
  assign T2692 = RouterBuffer_1_io_deq_bits_x[5'h1f:1'h1];
  assign T2693 = T2695 & T2694;
  assign T2694 = 3'h3 <= VCRouterStateManagement_1_io_currentState;
  assign T2695 = T2696;
  assign T2696 = R2697[1'h0:1'h0];
  assign T3186 = reset ? 8'h0 : T2698;
  assign T2698 = 1'h1 << CMeshDOR_1_io_result;
  assign T2699 = T2701 & T2700;
  assign T2700 = VCRouterStateManagement_1_io_currentState == 3'h4;
  assign T2701 = R2702;
  assign T3187 = reset ? 1'h1 : T1548;
  assign T3188 = reset ? 3'h0 : T2704;
  assign T2704 = T1382 ? T2705 : R2703;
  assign T2705 = T2706[2'h2:1'h0];
  assign T2706 = RouterBuffer_2_io_deq_bits_x[5'h1f:1'h1];
  assign T2707 = T2709 & T2708;
  assign T2708 = 3'h3 <= VCRouterStateManagement_2_io_currentState;
  assign T2709 = T2710;
  assign T2710 = R2711[1'h0:1'h0];
  assign T3189 = reset ? 8'h0 : T2712;
  assign T2712 = 1'h1 << CMeshDOR_2_io_result;
  assign T2713 = T2715 & T2714;
  assign T2714 = VCRouterStateManagement_2_io_currentState == 3'h4;
  assign T2715 = R2716;
  assign T3190 = reset ? 1'h1 : T1404;
  assign T3191 = reset ? 3'h0 : T2718;
  assign T2718 = T1238 ? T2719 : R2717;
  assign T2719 = T2720[2'h2:1'h0];
  assign T2720 = RouterBuffer_3_io_deq_bits_x[5'h1f:1'h1];
  assign T2721 = T2723 & T2722;
  assign T2722 = 3'h3 <= VCRouterStateManagement_3_io_currentState;
  assign T2723 = T2724;
  assign T2724 = R2725[1'h0:1'h0];
  assign T3192 = reset ? 8'h0 : T2726;
  assign T2726 = 1'h1 << CMeshDOR_3_io_result;
  assign T2727 = T2729 & T2728;
  assign T2728 = VCRouterStateManagement_3_io_currentState == 3'h4;
  assign T2729 = R2730;
  assign T3193 = reset ? 1'h1 : T1260;
  assign T3194 = reset ? 3'h0 : T2732;
  assign T2732 = T1094 ? T2733 : R2731;
  assign T2733 = T2734[2'h2:1'h0];
  assign T2734 = RouterBuffer_4_io_deq_bits_x[5'h1f:1'h1];
  assign T2735 = T2737 & T2736;
  assign T2736 = 3'h3 <= VCRouterStateManagement_4_io_currentState;
  assign T2737 = T2738;
  assign T2738 = R2739[1'h0:1'h0];
  assign T3195 = reset ? 8'h0 : T2740;
  assign T2740 = 1'h1 << CMeshDOR_4_io_result;
  assign T2741 = T2743 & T2742;
  assign T2742 = VCRouterStateManagement_4_io_currentState == 3'h4;
  assign T2743 = R2744;
  assign T3196 = reset ? 1'h1 : T1116;
  assign T3197 = reset ? 3'h0 : T2746;
  assign T2746 = T950 ? T2747 : R2745;
  assign T2747 = T2748[2'h2:1'h0];
  assign T2748 = RouterBuffer_5_io_deq_bits_x[5'h1f:1'h1];
  assign T2749 = T2751 & T2750;
  assign T2750 = 3'h3 <= VCRouterStateManagement_5_io_currentState;
  assign T2751 = T2752;
  assign T2752 = R2753[1'h0:1'h0];
  assign T3198 = reset ? 8'h0 : T2754;
  assign T2754 = 1'h1 << CMeshDOR_5_io_result;
  assign T2755 = T2757 & T2756;
  assign T2756 = VCRouterStateManagement_5_io_currentState == 3'h4;
  assign T2757 = R2758;
  assign T3199 = reset ? 1'h1 : T972;
  assign T3200 = reset ? 3'h0 : T2760;
  assign T2760 = T806 ? T2761 : R2759;
  assign T2761 = T2762[2'h2:1'h0];
  assign T2762 = RouterBuffer_6_io_deq_bits_x[5'h1f:1'h1];
  assign T2763 = T2765 & T2764;
  assign T2764 = 3'h3 <= VCRouterStateManagement_6_io_currentState;
  assign T2765 = T2766;
  assign T2766 = R2767[1'h0:1'h0];
  assign T3201 = reset ? 8'h0 : T2768;
  assign T2768 = 1'h1 << CMeshDOR_6_io_result;
  assign T2769 = T2771 & T2770;
  assign T2770 = VCRouterStateManagement_6_io_currentState == 3'h4;
  assign T2771 = R2772;
  assign T3202 = reset ? 1'h1 : T828;
  assign T3203 = reset ? 3'h0 : T2774;
  assign T2774 = T662 ? T2775 : R2773;
  assign T2775 = T2776[2'h2:1'h0];
  assign T2776 = RouterBuffer_7_io_deq_bits_x[5'h1f:1'h1];
  assign T2777 = T2779 & T2778;
  assign T2778 = 3'h3 <= VCRouterStateManagement_7_io_currentState;
  assign T2779 = T2780;
  assign T2780 = R2781[1'h0:1'h0];
  assign T3204 = reset ? 8'h0 : T2782;
  assign T2782 = 1'h1 << CMeshDOR_7_io_result;
  assign T2783 = T2785 & T2784;
  assign T2784 = VCRouterStateManagement_7_io_currentState == 3'h4;
  assign T2785 = R2786;
  assign T3205 = reset ? 1'h1 : T684;
  assign T3206 = reset ? 3'h0 : T2788;
  assign T2788 = T518 ? T2789 : R2787;
  assign T2789 = T2790[2'h2:1'h0];
  assign T2790 = RouterBuffer_8_io_deq_bits_x[5'h1f:1'h1];
  assign T2791 = T2793 & T2792;
  assign T2792 = 3'h3 <= VCRouterStateManagement_8_io_currentState;
  assign T2793 = T2794;
  assign T2794 = R2795[1'h0:1'h0];
  assign T3207 = reset ? 8'h0 : T2796;
  assign T2796 = 1'h1 << CMeshDOR_8_io_result;
  assign T2797 = T2799 & T2798;
  assign T2798 = VCRouterStateManagement_8_io_currentState == 3'h4;
  assign T2799 = R2800;
  assign T3208 = reset ? 1'h1 : T540;
  assign T3209 = reset ? 3'h0 : T2802;
  assign T2802 = T374 ? T2803 : R2801;
  assign T2803 = T2804[2'h2:1'h0];
  assign T2804 = RouterBuffer_9_io_deq_bits_x[5'h1f:1'h1];
  assign T2805 = T2807 & T2806;
  assign T2806 = 3'h3 <= VCRouterStateManagement_9_io_currentState;
  assign T2807 = T2808;
  assign T2808 = R2809[1'h0:1'h0];
  assign T3210 = reset ? 8'h0 : T2810;
  assign T2810 = 1'h1 << CMeshDOR_9_io_result;
  assign T2811 = T2813 & T2812;
  assign T2812 = VCRouterStateManagement_9_io_currentState == 3'h4;
  assign T2813 = R2814;
  assign T3211 = reset ? 1'h1 : T396;
  assign T2815 = T2817 & T2816;
  assign T2816 = 3'h3 <= VCRouterStateManagement_io_currentState;
  assign T2817 = T2818;
  assign T2818 = R2683[1'h1:1'h1];
  assign T2819 = T2821 & T2820;
  assign T2820 = VCRouterStateManagement_io_currentState == 3'h4;
  assign T2821 = R2688;
  assign T2822 = T2824 & T2823;
  assign T2823 = 3'h3 <= VCRouterStateManagement_1_io_currentState;
  assign T2824 = T2825;
  assign T2825 = R2697[1'h1:1'h1];
  assign T2826 = T2828 & T2827;
  assign T2827 = VCRouterStateManagement_1_io_currentState == 3'h4;
  assign T2828 = R2702;
  assign T2829 = T2831 & T2830;
  assign T2830 = 3'h3 <= VCRouterStateManagement_2_io_currentState;
  assign T2831 = T2832;
  assign T2832 = R2711[1'h1:1'h1];
  assign T2833 = T2835 & T2834;
  assign T2834 = VCRouterStateManagement_2_io_currentState == 3'h4;
  assign T2835 = R2716;
  assign T2836 = T2838 & T2837;
  assign T2837 = 3'h3 <= VCRouterStateManagement_3_io_currentState;
  assign T2838 = T2839;
  assign T2839 = R2725[1'h1:1'h1];
  assign T2840 = T2842 & T2841;
  assign T2841 = VCRouterStateManagement_3_io_currentState == 3'h4;
  assign T2842 = R2730;
  assign T2843 = T2845 & T2844;
  assign T2844 = 3'h3 <= VCRouterStateManagement_4_io_currentState;
  assign T2845 = T2846;
  assign T2846 = R2739[1'h1:1'h1];
  assign T2847 = T2849 & T2848;
  assign T2848 = VCRouterStateManagement_4_io_currentState == 3'h4;
  assign T2849 = R2744;
  assign T2850 = T2852 & T2851;
  assign T2851 = 3'h3 <= VCRouterStateManagement_5_io_currentState;
  assign T2852 = T2853;
  assign T2853 = R2753[1'h1:1'h1];
  assign T2854 = T2856 & T2855;
  assign T2855 = VCRouterStateManagement_5_io_currentState == 3'h4;
  assign T2856 = R2758;
  assign T2857 = T2859 & T2858;
  assign T2858 = 3'h3 <= VCRouterStateManagement_6_io_currentState;
  assign T2859 = T2860;
  assign T2860 = R2767[1'h1:1'h1];
  assign T2861 = T2863 & T2862;
  assign T2862 = VCRouterStateManagement_6_io_currentState == 3'h4;
  assign T2863 = R2772;
  assign T2864 = T2866 & T2865;
  assign T2865 = 3'h3 <= VCRouterStateManagement_7_io_currentState;
  assign T2866 = T2867;
  assign T2867 = R2781[1'h1:1'h1];
  assign T2868 = T2870 & T2869;
  assign T2869 = VCRouterStateManagement_7_io_currentState == 3'h4;
  assign T2870 = R2786;
  assign T2871 = T2873 & T2872;
  assign T2872 = 3'h3 <= VCRouterStateManagement_8_io_currentState;
  assign T2873 = T2874;
  assign T2874 = R2795[1'h1:1'h1];
  assign T2875 = T2877 & T2876;
  assign T2876 = VCRouterStateManagement_8_io_currentState == 3'h4;
  assign T2877 = R2800;
  assign T2878 = T2880 & T2879;
  assign T2879 = 3'h3 <= VCRouterStateManagement_9_io_currentState;
  assign T2880 = T2881;
  assign T2881 = R2809[1'h1:1'h1];
  assign T2882 = T2884 & T2883;
  assign T2883 = VCRouterStateManagement_9_io_currentState == 3'h4;
  assign T2884 = R2814;
  assign T2885 = T2887 & T2886;
  assign T2886 = 3'h3 <= VCRouterStateManagement_io_currentState;
  assign T2887 = T2888;
  assign T2888 = R2683[2'h2:2'h2];
  assign T2889 = T2891 & T2890;
  assign T2890 = VCRouterStateManagement_io_currentState == 3'h4;
  assign T2891 = R2688;
  assign T2892 = T2894 & T2893;
  assign T2893 = 3'h3 <= VCRouterStateManagement_1_io_currentState;
  assign T2894 = T2895;
  assign T2895 = R2697[2'h2:2'h2];
  assign T2896 = T2898 & T2897;
  assign T2897 = VCRouterStateManagement_1_io_currentState == 3'h4;
  assign T2898 = R2702;
  assign T2899 = T2901 & T2900;
  assign T2900 = 3'h3 <= VCRouterStateManagement_2_io_currentState;
  assign T2901 = T2902;
  assign T2902 = R2711[2'h2:2'h2];
  assign T2903 = T2905 & T2904;
  assign T2904 = VCRouterStateManagement_2_io_currentState == 3'h4;
  assign T2905 = R2716;
  assign T2906 = T2908 & T2907;
  assign T2907 = 3'h3 <= VCRouterStateManagement_3_io_currentState;
  assign T2908 = T2909;
  assign T2909 = R2725[2'h2:2'h2];
  assign T2910 = T2912 & T2911;
  assign T2911 = VCRouterStateManagement_3_io_currentState == 3'h4;
  assign T2912 = R2730;
  assign T2913 = T2915 & T2914;
  assign T2914 = 3'h3 <= VCRouterStateManagement_4_io_currentState;
  assign T2915 = T2916;
  assign T2916 = R2739[2'h2:2'h2];
  assign T2917 = T2919 & T2918;
  assign T2918 = VCRouterStateManagement_4_io_currentState == 3'h4;
  assign T2919 = R2744;
  assign T2920 = T2922 & T2921;
  assign T2921 = 3'h3 <= VCRouterStateManagement_5_io_currentState;
  assign T2922 = T2923;
  assign T2923 = R2753[2'h2:2'h2];
  assign T2924 = T2926 & T2925;
  assign T2925 = VCRouterStateManagement_5_io_currentState == 3'h4;
  assign T2926 = R2758;
  assign T2927 = T2929 & T2928;
  assign T2928 = 3'h3 <= VCRouterStateManagement_6_io_currentState;
  assign T2929 = T2930;
  assign T2930 = R2767[2'h2:2'h2];
  assign T2931 = T2933 & T2932;
  assign T2932 = VCRouterStateManagement_6_io_currentState == 3'h4;
  assign T2933 = R2772;
  assign T2934 = T2936 & T2935;
  assign T2935 = 3'h3 <= VCRouterStateManagement_7_io_currentState;
  assign T2936 = T2937;
  assign T2937 = R2781[2'h2:2'h2];
  assign T2938 = T2940 & T2939;
  assign T2939 = VCRouterStateManagement_7_io_currentState == 3'h4;
  assign T2940 = R2786;
  assign T2941 = T2943 & T2942;
  assign T2942 = 3'h3 <= VCRouterStateManagement_8_io_currentState;
  assign T2943 = T2944;
  assign T2944 = R2795[2'h2:2'h2];
  assign T2945 = T2947 & T2946;
  assign T2946 = VCRouterStateManagement_8_io_currentState == 3'h4;
  assign T2947 = R2800;
  assign T2948 = T2950 & T2949;
  assign T2949 = 3'h3 <= VCRouterStateManagement_9_io_currentState;
  assign T2950 = T2951;
  assign T2951 = R2809[2'h2:2'h2];
  assign T2952 = T2954 & T2953;
  assign T2953 = VCRouterStateManagement_9_io_currentState == 3'h4;
  assign T2954 = R2814;
  assign T2955 = T2957 & T2956;
  assign T2956 = 3'h3 <= VCRouterStateManagement_io_currentState;
  assign T2957 = T2958;
  assign T2958 = R2683[2'h3:2'h3];
  assign T2959 = T2961 & T2960;
  assign T2960 = VCRouterStateManagement_io_currentState == 3'h4;
  assign T2961 = R2688;
  assign T2962 = T2964 & T2963;
  assign T2963 = 3'h3 <= VCRouterStateManagement_1_io_currentState;
  assign T2964 = T2965;
  assign T2965 = R2697[2'h3:2'h3];
  assign T2966 = T2968 & T2967;
  assign T2967 = VCRouterStateManagement_1_io_currentState == 3'h4;
  assign T2968 = R2702;
  assign T2969 = T2971 & T2970;
  assign T2970 = 3'h3 <= VCRouterStateManagement_2_io_currentState;
  assign T2971 = T2972;
  assign T2972 = R2711[2'h3:2'h3];
  assign T2973 = T2975 & T2974;
  assign T2974 = VCRouterStateManagement_2_io_currentState == 3'h4;
  assign T2975 = R2716;
  assign T2976 = T2978 & T2977;
  assign T2977 = 3'h3 <= VCRouterStateManagement_3_io_currentState;
  assign T2978 = T2979;
  assign T2979 = R2725[2'h3:2'h3];
  assign T2980 = T2982 & T2981;
  assign T2981 = VCRouterStateManagement_3_io_currentState == 3'h4;
  assign T2982 = R2730;
  assign T2983 = T2985 & T2984;
  assign T2984 = 3'h3 <= VCRouterStateManagement_4_io_currentState;
  assign T2985 = T2986;
  assign T2986 = R2739[2'h3:2'h3];
  assign T2987 = T2989 & T2988;
  assign T2988 = VCRouterStateManagement_4_io_currentState == 3'h4;
  assign T2989 = R2744;
  assign T2990 = T2992 & T2991;
  assign T2991 = 3'h3 <= VCRouterStateManagement_5_io_currentState;
  assign T2992 = T2993;
  assign T2993 = R2753[2'h3:2'h3];
  assign T2994 = T2996 & T2995;
  assign T2995 = VCRouterStateManagement_5_io_currentState == 3'h4;
  assign T2996 = R2758;
  assign T2997 = T2999 & T2998;
  assign T2998 = 3'h3 <= VCRouterStateManagement_6_io_currentState;
  assign T2999 = T3000;
  assign T3000 = R2767[2'h3:2'h3];
  assign T3001 = T3003 & T3002;
  assign T3002 = VCRouterStateManagement_6_io_currentState == 3'h4;
  assign T3003 = R2772;
  assign T3004 = T3006 & T3005;
  assign T3005 = 3'h3 <= VCRouterStateManagement_7_io_currentState;
  assign T3006 = T3007;
  assign T3007 = R2781[2'h3:2'h3];
  assign T3008 = T3010 & T3009;
  assign T3009 = VCRouterStateManagement_7_io_currentState == 3'h4;
  assign T3010 = R2786;
  assign T3011 = T3013 & T3012;
  assign T3012 = 3'h3 <= VCRouterStateManagement_8_io_currentState;
  assign T3013 = T3014;
  assign T3014 = R2795[2'h3:2'h3];
  assign T3015 = T3017 & T3016;
  assign T3016 = VCRouterStateManagement_8_io_currentState == 3'h4;
  assign T3017 = R2800;
  assign T3018 = T3020 & T3019;
  assign T3019 = 3'h3 <= VCRouterStateManagement_9_io_currentState;
  assign T3020 = T3021;
  assign T3021 = R2809[2'h3:2'h3];
  assign T3022 = T3024 & T3023;
  assign T3023 = VCRouterStateManagement_9_io_currentState == 3'h4;
  assign T3024 = R2814;
  assign T3025 = T3027 & T3026;
  assign T3026 = 3'h3 <= VCRouterStateManagement_io_currentState;
  assign T3027 = T3028;
  assign T3028 = R2683[3'h4:3'h4];
  assign T3029 = T3031 & T3030;
  assign T3030 = VCRouterStateManagement_io_currentState == 3'h4;
  assign T3031 = R2688;
  assign T3032 = T3034 & T3033;
  assign T3033 = 3'h3 <= VCRouterStateManagement_1_io_currentState;
  assign T3034 = T3035;
  assign T3035 = R2697[3'h4:3'h4];
  assign T3036 = T3038 & T3037;
  assign T3037 = VCRouterStateManagement_1_io_currentState == 3'h4;
  assign T3038 = R2702;
  assign T3039 = T3041 & T3040;
  assign T3040 = 3'h3 <= VCRouterStateManagement_2_io_currentState;
  assign T3041 = T3042;
  assign T3042 = R2711[3'h4:3'h4];
  assign T3043 = T3045 & T3044;
  assign T3044 = VCRouterStateManagement_2_io_currentState == 3'h4;
  assign T3045 = R2716;
  assign T3046 = T3048 & T3047;
  assign T3047 = 3'h3 <= VCRouterStateManagement_3_io_currentState;
  assign T3048 = T3049;
  assign T3049 = R2725[3'h4:3'h4];
  assign T3050 = T3052 & T3051;
  assign T3051 = VCRouterStateManagement_3_io_currentState == 3'h4;
  assign T3052 = R2730;
  assign T3053 = T3055 & T3054;
  assign T3054 = 3'h3 <= VCRouterStateManagement_4_io_currentState;
  assign T3055 = T3056;
  assign T3056 = R2739[3'h4:3'h4];
  assign T3057 = T3059 & T3058;
  assign T3058 = VCRouterStateManagement_4_io_currentState == 3'h4;
  assign T3059 = R2744;
  assign T3060 = T3062 & T3061;
  assign T3061 = 3'h3 <= VCRouterStateManagement_5_io_currentState;
  assign T3062 = T3063;
  assign T3063 = R2753[3'h4:3'h4];
  assign T3064 = T3066 & T3065;
  assign T3065 = VCRouterStateManagement_5_io_currentState == 3'h4;
  assign T3066 = R2758;
  assign T3067 = T3069 & T3068;
  assign T3068 = 3'h3 <= VCRouterStateManagement_6_io_currentState;
  assign T3069 = T3070;
  assign T3070 = R2767[3'h4:3'h4];
  assign T3071 = T3073 & T3072;
  assign T3072 = VCRouterStateManagement_6_io_currentState == 3'h4;
  assign T3073 = R2772;
  assign T3074 = T3076 & T3075;
  assign T3075 = 3'h3 <= VCRouterStateManagement_7_io_currentState;
  assign T3076 = T3077;
  assign T3077 = R2781[3'h4:3'h4];
  assign T3078 = T3080 & T3079;
  assign T3079 = VCRouterStateManagement_7_io_currentState == 3'h4;
  assign T3080 = R2786;
  assign T3081 = T3083 & T3082;
  assign T3082 = 3'h3 <= VCRouterStateManagement_8_io_currentState;
  assign T3083 = T3084;
  assign T3084 = R2795[3'h4:3'h4];
  assign T3085 = T3087 & T3086;
  assign T3086 = VCRouterStateManagement_8_io_currentState == 3'h4;
  assign T3087 = R2800;
  assign T3088 = T3090 & T3089;
  assign T3089 = 3'h3 <= VCRouterStateManagement_9_io_currentState;
  assign T3090 = T3091;
  assign T3091 = R2809[3'h4:3'h4];
  assign T3092 = T3094 & T3093;
  assign T3093 = VCRouterStateManagement_9_io_currentState == 3'h4;
  assign T3094 = R2814;
  assign io_counters_0_counterVal = T3212;
  assign T3212 = {31'h0, T3095};
  assign T3095 = T3096 == 1'h0;
  assign T3096 = T365 ^ 1'h1;
  assign io_outChannels_0_flitValid = R3097;
  assign io_outChannels_0_flit_x = R3098;
  assign T3099 = 55'h0;
  assign T3213 = reset ? T3099 : switch_io_outPorts_0_x;
  assign io_outChannels_1_flitValid = R3100;
  assign io_outChannels_1_flit_x = R3101;
  assign T3102 = 55'h0;
  assign T3214 = reset ? T3102 : switch_io_outPorts_1_x;
  assign io_outChannels_2_flitValid = R3103;
  assign io_outChannels_2_flit_x = R3104;
  assign T3105 = 55'h0;
  assign T3215 = reset ? T3105 : switch_io_outPorts_2_x;
  assign io_outChannels_3_flitValid = R3106;
  assign io_outChannels_3_flit_x = R3107;
  assign T3108 = 55'h0;
  assign T3216 = reset ? T3108 : switch_io_outPorts_3_x;
  assign io_outChannels_4_flitValid = R3109;
  assign io_outChannels_4_flit_x = R3110;
  assign T3111 = 55'h0;
  assign T3217 = reset ? T3111 : switch_io_outPorts_4_x;
  assign io_inChannels_0_credit_0_grant = CreditGen_io_outCredit_grant;
  assign io_inChannels_0_credit_1_grant = CreditGen_1_io_outCredit_grant;
  assign io_inChannels_1_credit_0_grant = CreditGen_2_io_outCredit_grant;
  assign io_inChannels_1_credit_1_grant = CreditGen_3_io_outCredit_grant;
  assign io_inChannels_2_credit_0_grant = CreditGen_4_io_outCredit_grant;
  assign io_inChannels_2_credit_1_grant = CreditGen_5_io_outCredit_grant;
  assign io_inChannels_3_credit_0_grant = CreditGen_6_io_outCredit_grant;
  assign io_inChannels_3_credit_1_grant = CreditGen_7_io_outCredit_grant;
  assign io_inChannels_4_credit_0_grant = CreditGen_8_io_outCredit_grant;
  assign io_inChannels_4_credit_1_grant = CreditGen_9_io_outCredit_grant;
  Switch switch(
       .io_inPorts_9_x( ReplaceVCPort_9_io_newFlit_x ),
       .io_inPorts_8_x( ReplaceVCPort_8_io_newFlit_x ),
       .io_inPorts_7_x( ReplaceVCPort_7_io_newFlit_x ),
       .io_inPorts_6_x( ReplaceVCPort_6_io_newFlit_x ),
       .io_inPorts_5_x( ReplaceVCPort_5_io_newFlit_x ),
       .io_inPorts_4_x( ReplaceVCPort_4_io_newFlit_x ),
       .io_inPorts_3_x( ReplaceVCPort_3_io_newFlit_x ),
       .io_inPorts_2_x( ReplaceVCPort_2_io_newFlit_x ),
       .io_inPorts_1_x( ReplaceVCPort_1_io_newFlit_x ),
       .io_inPorts_0_x( ReplaceVCPort_io_newFlit_x ),
       .io_outPorts_4_x( switch_io_outPorts_4_x ),
       .io_outPorts_3_x( switch_io_outPorts_3_x ),
       .io_outPorts_2_x( switch_io_outPorts_2_x ),
       .io_outPorts_1_x( switch_io_outPorts_1_x ),
       .io_outPorts_0_x( switch_io_outPorts_0_x ),
       .io_sel_4( swAllocator_io_chosens_4 ),
       .io_sel_3( swAllocator_io_chosens_3 ),
       .io_sel_2( swAllocator_io_chosens_2 ),
       .io_sel_1( swAllocator_io_chosens_1 ),
       .io_sel_0( swAllocator_io_chosens_0 )
  );
  SwitchAllocator_0 swAllocator(.clk(clk), .reset(reset),
       .io_requests_4_9_releaseLock( T3092 ),
       .io_requests_4_9_grant( swAllocator_io_requests_4_9_grant ),
       .io_requests_4_9_request( T3088 ),
       .io_requests_4_9_priorityLevel( R2801 ),
       .io_requests_4_8_releaseLock( T3085 ),
       .io_requests_4_8_grant( swAllocator_io_requests_4_8_grant ),
       .io_requests_4_8_request( T3081 ),
       .io_requests_4_8_priorityLevel( R2787 ),
       .io_requests_4_7_releaseLock( T3078 ),
       .io_requests_4_7_grant( swAllocator_io_requests_4_7_grant ),
       .io_requests_4_7_request( T3074 ),
       .io_requests_4_7_priorityLevel( R2773 ),
       .io_requests_4_6_releaseLock( T3071 ),
       .io_requests_4_6_grant( swAllocator_io_requests_4_6_grant ),
       .io_requests_4_6_request( T3067 ),
       .io_requests_4_6_priorityLevel( R2759 ),
       .io_requests_4_5_releaseLock( T3064 ),
       .io_requests_4_5_grant( swAllocator_io_requests_4_5_grant ),
       .io_requests_4_5_request( T3060 ),
       .io_requests_4_5_priorityLevel( R2745 ),
       .io_requests_4_4_releaseLock( T3057 ),
       .io_requests_4_4_grant( swAllocator_io_requests_4_4_grant ),
       .io_requests_4_4_request( T3053 ),
       .io_requests_4_4_priorityLevel( R2731 ),
       .io_requests_4_3_releaseLock( T3050 ),
       .io_requests_4_3_grant( swAllocator_io_requests_4_3_grant ),
       .io_requests_4_3_request( T3046 ),
       .io_requests_4_3_priorityLevel( R2717 ),
       .io_requests_4_2_releaseLock( T3043 ),
       .io_requests_4_2_grant( swAllocator_io_requests_4_2_grant ),
       .io_requests_4_2_request( T3039 ),
       .io_requests_4_2_priorityLevel( R2703 ),
       .io_requests_4_1_releaseLock( T3036 ),
       .io_requests_4_1_grant( swAllocator_io_requests_4_1_grant ),
       .io_requests_4_1_request( T3032 ),
       .io_requests_4_1_priorityLevel( R2689 ),
       .io_requests_4_0_releaseLock( T3029 ),
       .io_requests_4_0_grant( swAllocator_io_requests_4_0_grant ),
       .io_requests_4_0_request( T3025 ),
       .io_requests_4_0_priorityLevel( R2675 ),
       .io_requests_3_9_releaseLock( T3022 ),
       .io_requests_3_9_grant( swAllocator_io_requests_3_9_grant ),
       .io_requests_3_9_request( T3018 ),
       .io_requests_3_9_priorityLevel( R2801 ),
       .io_requests_3_8_releaseLock( T3015 ),
       .io_requests_3_8_grant( swAllocator_io_requests_3_8_grant ),
       .io_requests_3_8_request( T3011 ),
       .io_requests_3_8_priorityLevel( R2787 ),
       .io_requests_3_7_releaseLock( T3008 ),
       .io_requests_3_7_grant( swAllocator_io_requests_3_7_grant ),
       .io_requests_3_7_request( T3004 ),
       .io_requests_3_7_priorityLevel( R2773 ),
       .io_requests_3_6_releaseLock( T3001 ),
       .io_requests_3_6_grant( swAllocator_io_requests_3_6_grant ),
       .io_requests_3_6_request( T2997 ),
       .io_requests_3_6_priorityLevel( R2759 ),
       .io_requests_3_5_releaseLock( T2994 ),
       .io_requests_3_5_grant( swAllocator_io_requests_3_5_grant ),
       .io_requests_3_5_request( T2990 ),
       .io_requests_3_5_priorityLevel( R2745 ),
       .io_requests_3_4_releaseLock( T2987 ),
       .io_requests_3_4_grant( swAllocator_io_requests_3_4_grant ),
       .io_requests_3_4_request( T2983 ),
       .io_requests_3_4_priorityLevel( R2731 ),
       .io_requests_3_3_releaseLock( T2980 ),
       .io_requests_3_3_grant( swAllocator_io_requests_3_3_grant ),
       .io_requests_3_3_request( T2976 ),
       .io_requests_3_3_priorityLevel( R2717 ),
       .io_requests_3_2_releaseLock( T2973 ),
       .io_requests_3_2_grant( swAllocator_io_requests_3_2_grant ),
       .io_requests_3_2_request( T2969 ),
       .io_requests_3_2_priorityLevel( R2703 ),
       .io_requests_3_1_releaseLock( T2966 ),
       .io_requests_3_1_grant( swAllocator_io_requests_3_1_grant ),
       .io_requests_3_1_request( T2962 ),
       .io_requests_3_1_priorityLevel( R2689 ),
       .io_requests_3_0_releaseLock( T2959 ),
       .io_requests_3_0_grant( swAllocator_io_requests_3_0_grant ),
       .io_requests_3_0_request( T2955 ),
       .io_requests_3_0_priorityLevel( R2675 ),
       .io_requests_2_9_releaseLock( T2952 ),
       .io_requests_2_9_grant( swAllocator_io_requests_2_9_grant ),
       .io_requests_2_9_request( T2948 ),
       .io_requests_2_9_priorityLevel( R2801 ),
       .io_requests_2_8_releaseLock( T2945 ),
       .io_requests_2_8_grant( swAllocator_io_requests_2_8_grant ),
       .io_requests_2_8_request( T2941 ),
       .io_requests_2_8_priorityLevel( R2787 ),
       .io_requests_2_7_releaseLock( T2938 ),
       .io_requests_2_7_grant( swAllocator_io_requests_2_7_grant ),
       .io_requests_2_7_request( T2934 ),
       .io_requests_2_7_priorityLevel( R2773 ),
       .io_requests_2_6_releaseLock( T2931 ),
       .io_requests_2_6_grant( swAllocator_io_requests_2_6_grant ),
       .io_requests_2_6_request( T2927 ),
       .io_requests_2_6_priorityLevel( R2759 ),
       .io_requests_2_5_releaseLock( T2924 ),
       .io_requests_2_5_grant( swAllocator_io_requests_2_5_grant ),
       .io_requests_2_5_request( T2920 ),
       .io_requests_2_5_priorityLevel( R2745 ),
       .io_requests_2_4_releaseLock( T2917 ),
       .io_requests_2_4_grant( swAllocator_io_requests_2_4_grant ),
       .io_requests_2_4_request( T2913 ),
       .io_requests_2_4_priorityLevel( R2731 ),
       .io_requests_2_3_releaseLock( T2910 ),
       .io_requests_2_3_grant( swAllocator_io_requests_2_3_grant ),
       .io_requests_2_3_request( T2906 ),
       .io_requests_2_3_priorityLevel( R2717 ),
       .io_requests_2_2_releaseLock( T2903 ),
       .io_requests_2_2_grant( swAllocator_io_requests_2_2_grant ),
       .io_requests_2_2_request( T2899 ),
       .io_requests_2_2_priorityLevel( R2703 ),
       .io_requests_2_1_releaseLock( T2896 ),
       .io_requests_2_1_grant( swAllocator_io_requests_2_1_grant ),
       .io_requests_2_1_request( T2892 ),
       .io_requests_2_1_priorityLevel( R2689 ),
       .io_requests_2_0_releaseLock( T2889 ),
       .io_requests_2_0_grant( swAllocator_io_requests_2_0_grant ),
       .io_requests_2_0_request( T2885 ),
       .io_requests_2_0_priorityLevel( R2675 ),
       .io_requests_1_9_releaseLock( T2882 ),
       .io_requests_1_9_grant( swAllocator_io_requests_1_9_grant ),
       .io_requests_1_9_request( T2878 ),
       .io_requests_1_9_priorityLevel( R2801 ),
       .io_requests_1_8_releaseLock( T2875 ),
       .io_requests_1_8_grant( swAllocator_io_requests_1_8_grant ),
       .io_requests_1_8_request( T2871 ),
       .io_requests_1_8_priorityLevel( R2787 ),
       .io_requests_1_7_releaseLock( T2868 ),
       .io_requests_1_7_grant( swAllocator_io_requests_1_7_grant ),
       .io_requests_1_7_request( T2864 ),
       .io_requests_1_7_priorityLevel( R2773 ),
       .io_requests_1_6_releaseLock( T2861 ),
       .io_requests_1_6_grant( swAllocator_io_requests_1_6_grant ),
       .io_requests_1_6_request( T2857 ),
       .io_requests_1_6_priorityLevel( R2759 ),
       .io_requests_1_5_releaseLock( T2854 ),
       .io_requests_1_5_grant( swAllocator_io_requests_1_5_grant ),
       .io_requests_1_5_request( T2850 ),
       .io_requests_1_5_priorityLevel( R2745 ),
       .io_requests_1_4_releaseLock( T2847 ),
       .io_requests_1_4_grant( swAllocator_io_requests_1_4_grant ),
       .io_requests_1_4_request( T2843 ),
       .io_requests_1_4_priorityLevel( R2731 ),
       .io_requests_1_3_releaseLock( T2840 ),
       .io_requests_1_3_grant( swAllocator_io_requests_1_3_grant ),
       .io_requests_1_3_request( T2836 ),
       .io_requests_1_3_priorityLevel( R2717 ),
       .io_requests_1_2_releaseLock( T2833 ),
       .io_requests_1_2_grant( swAllocator_io_requests_1_2_grant ),
       .io_requests_1_2_request( T2829 ),
       .io_requests_1_2_priorityLevel( R2703 ),
       .io_requests_1_1_releaseLock( T2826 ),
       .io_requests_1_1_grant( swAllocator_io_requests_1_1_grant ),
       .io_requests_1_1_request( T2822 ),
       .io_requests_1_1_priorityLevel( R2689 ),
       .io_requests_1_0_releaseLock( T2819 ),
       .io_requests_1_0_grant( swAllocator_io_requests_1_0_grant ),
       .io_requests_1_0_request( T2815 ),
       .io_requests_1_0_priorityLevel( R2675 ),
       .io_requests_0_9_releaseLock( T2811 ),
       .io_requests_0_9_grant( swAllocator_io_requests_0_9_grant ),
       .io_requests_0_9_request( T2805 ),
       .io_requests_0_9_priorityLevel( R2801 ),
       .io_requests_0_8_releaseLock( T2797 ),
       .io_requests_0_8_grant( swAllocator_io_requests_0_8_grant ),
       .io_requests_0_8_request( T2791 ),
       .io_requests_0_8_priorityLevel( R2787 ),
       .io_requests_0_7_releaseLock( T2783 ),
       .io_requests_0_7_grant( swAllocator_io_requests_0_7_grant ),
       .io_requests_0_7_request( T2777 ),
       .io_requests_0_7_priorityLevel( R2773 ),
       .io_requests_0_6_releaseLock( T2769 ),
       .io_requests_0_6_grant( swAllocator_io_requests_0_6_grant ),
       .io_requests_0_6_request( T2763 ),
       .io_requests_0_6_priorityLevel( R2759 ),
       .io_requests_0_5_releaseLock( T2755 ),
       .io_requests_0_5_grant( swAllocator_io_requests_0_5_grant ),
       .io_requests_0_5_request( T2749 ),
       .io_requests_0_5_priorityLevel( R2745 ),
       .io_requests_0_4_releaseLock( T2741 ),
       .io_requests_0_4_grant( swAllocator_io_requests_0_4_grant ),
       .io_requests_0_4_request( T2735 ),
       .io_requests_0_4_priorityLevel( R2731 ),
       .io_requests_0_3_releaseLock( T2727 ),
       .io_requests_0_3_grant( swAllocator_io_requests_0_3_grant ),
       .io_requests_0_3_request( T2721 ),
       .io_requests_0_3_priorityLevel( R2717 ),
       .io_requests_0_2_releaseLock( T2713 ),
       .io_requests_0_2_grant( swAllocator_io_requests_0_2_grant ),
       .io_requests_0_2_request( T2707 ),
       .io_requests_0_2_priorityLevel( R2703 ),
       .io_requests_0_1_releaseLock( T2699 ),
       .io_requests_0_1_grant( swAllocator_io_requests_0_1_grant ),
       .io_requests_0_1_request( T2693 ),
       .io_requests_0_1_priorityLevel( R2689 ),
       .io_requests_0_0_releaseLock( T2685 ),
       .io_requests_0_0_grant( swAllocator_io_requests_0_0_grant ),
       .io_requests_0_0_request( T2679 ),
       .io_requests_0_0_priorityLevel( R2675 ),
       .io_resources_4_ready( 1'h1 ),
       //.io_resources_4_valid(  )
       .io_resources_3_ready( 1'h1 ),
       //.io_resources_3_valid(  )
       .io_resources_2_ready( 1'h1 ),
       //.io_resources_2_valid(  )
       .io_resources_1_ready( 1'h1 ),
       //.io_resources_1_valid(  )
       .io_resources_0_ready( 1'h1 ),
       //.io_resources_0_valid(  )
       .io_chosens_4( swAllocator_io_chosens_4 ),
       .io_chosens_3( swAllocator_io_chosens_3 ),
       .io_chosens_2( swAllocator_io_chosens_2 ),
       .io_chosens_1( swAllocator_io_chosens_1 ),
       .io_chosens_0( swAllocator_io_chosens_0 )
  );
  SwitchAllocator_1 vcAllocator(.clk(clk), .reset(reset),
       .io_requests_9_9_releaseLock( R2671 ),
       //.io_requests_9_9_grant(  )
       .io_requests_9_9_request( T2670 ),
       //.io_requests_9_9_priorityLevel(  )
       .io_requests_9_8_releaseLock( R2666 ),
       //.io_requests_9_8_grant(  )
       .io_requests_9_8_request( T2665 ),
       //.io_requests_9_8_priorityLevel(  )
       .io_requests_9_7_releaseLock( R2661 ),
       //.io_requests_9_7_grant(  )
       .io_requests_9_7_request( T2660 ),
       //.io_requests_9_7_priorityLevel(  )
       .io_requests_9_6_releaseLock( R2656 ),
       //.io_requests_9_6_grant(  )
       .io_requests_9_6_request( T2655 ),
       //.io_requests_9_6_priorityLevel(  )
       .io_requests_9_5_releaseLock( R2651 ),
       //.io_requests_9_5_grant(  )
       .io_requests_9_5_request( T2650 ),
       //.io_requests_9_5_priorityLevel(  )
       .io_requests_9_4_releaseLock( R2646 ),
       //.io_requests_9_4_grant(  )
       .io_requests_9_4_request( T2645 ),
       //.io_requests_9_4_priorityLevel(  )
       .io_requests_9_3_releaseLock( R2641 ),
       //.io_requests_9_3_grant(  )
       .io_requests_9_3_request( T2640 ),
       //.io_requests_9_3_priorityLevel(  )
       .io_requests_9_2_releaseLock( R2636 ),
       //.io_requests_9_2_grant(  )
       .io_requests_9_2_request( T2635 ),
       //.io_requests_9_2_priorityLevel(  )
       .io_requests_9_1_releaseLock( R2631 ),
       //.io_requests_9_1_grant(  )
       .io_requests_9_1_request( T2630 ),
       //.io_requests_9_1_priorityLevel(  )
       .io_requests_9_0_releaseLock( R2626 ),
       //.io_requests_9_0_grant(  )
       .io_requests_9_0_request( T2625 ),
       //.io_requests_9_0_priorityLevel(  )
       .io_requests_8_9_releaseLock( R2621 ),
       //.io_requests_8_9_grant(  )
       .io_requests_8_9_request( T2620 ),
       //.io_requests_8_9_priorityLevel(  )
       .io_requests_8_8_releaseLock( R2616 ),
       //.io_requests_8_8_grant(  )
       .io_requests_8_8_request( T2615 ),
       //.io_requests_8_8_priorityLevel(  )
       .io_requests_8_7_releaseLock( R2611 ),
       //.io_requests_8_7_grant(  )
       .io_requests_8_7_request( T2610 ),
       //.io_requests_8_7_priorityLevel(  )
       .io_requests_8_6_releaseLock( R2606 ),
       //.io_requests_8_6_grant(  )
       .io_requests_8_6_request( T2605 ),
       //.io_requests_8_6_priorityLevel(  )
       .io_requests_8_5_releaseLock( R2601 ),
       //.io_requests_8_5_grant(  )
       .io_requests_8_5_request( T2600 ),
       //.io_requests_8_5_priorityLevel(  )
       .io_requests_8_4_releaseLock( R2596 ),
       //.io_requests_8_4_grant(  )
       .io_requests_8_4_request( T2595 ),
       //.io_requests_8_4_priorityLevel(  )
       .io_requests_8_3_releaseLock( R2591 ),
       //.io_requests_8_3_grant(  )
       .io_requests_8_3_request( T2590 ),
       //.io_requests_8_3_priorityLevel(  )
       .io_requests_8_2_releaseLock( R2586 ),
       //.io_requests_8_2_grant(  )
       .io_requests_8_2_request( T2585 ),
       //.io_requests_8_2_priorityLevel(  )
       .io_requests_8_1_releaseLock( R2581 ),
       //.io_requests_8_1_grant(  )
       .io_requests_8_1_request( T2580 ),
       //.io_requests_8_1_priorityLevel(  )
       .io_requests_8_0_releaseLock( R2576 ),
       //.io_requests_8_0_grant(  )
       .io_requests_8_0_request( T2575 ),
       //.io_requests_8_0_priorityLevel(  )
       .io_requests_7_9_releaseLock( R2571 ),
       //.io_requests_7_9_grant(  )
       .io_requests_7_9_request( T2570 ),
       //.io_requests_7_9_priorityLevel(  )
       .io_requests_7_8_releaseLock( R2566 ),
       //.io_requests_7_8_grant(  )
       .io_requests_7_8_request( T2565 ),
       //.io_requests_7_8_priorityLevel(  )
       .io_requests_7_7_releaseLock( R2561 ),
       //.io_requests_7_7_grant(  )
       .io_requests_7_7_request( T2560 ),
       //.io_requests_7_7_priorityLevel(  )
       .io_requests_7_6_releaseLock( R2556 ),
       //.io_requests_7_6_grant(  )
       .io_requests_7_6_request( T2555 ),
       //.io_requests_7_6_priorityLevel(  )
       .io_requests_7_5_releaseLock( R2551 ),
       //.io_requests_7_5_grant(  )
       .io_requests_7_5_request( T2550 ),
       //.io_requests_7_5_priorityLevel(  )
       .io_requests_7_4_releaseLock( R2546 ),
       //.io_requests_7_4_grant(  )
       .io_requests_7_4_request( T2545 ),
       //.io_requests_7_4_priorityLevel(  )
       .io_requests_7_3_releaseLock( R2541 ),
       //.io_requests_7_3_grant(  )
       .io_requests_7_3_request( T2540 ),
       //.io_requests_7_3_priorityLevel(  )
       .io_requests_7_2_releaseLock( R2536 ),
       //.io_requests_7_2_grant(  )
       .io_requests_7_2_request( T2535 ),
       //.io_requests_7_2_priorityLevel(  )
       .io_requests_7_1_releaseLock( R2531 ),
       //.io_requests_7_1_grant(  )
       .io_requests_7_1_request( T2530 ),
       //.io_requests_7_1_priorityLevel(  )
       .io_requests_7_0_releaseLock( R2526 ),
       //.io_requests_7_0_grant(  )
       .io_requests_7_0_request( T2525 ),
       //.io_requests_7_0_priorityLevel(  )
       .io_requests_6_9_releaseLock( R2521 ),
       //.io_requests_6_9_grant(  )
       .io_requests_6_9_request( T2520 ),
       //.io_requests_6_9_priorityLevel(  )
       .io_requests_6_8_releaseLock( R2516 ),
       //.io_requests_6_8_grant(  )
       .io_requests_6_8_request( T2515 ),
       //.io_requests_6_8_priorityLevel(  )
       .io_requests_6_7_releaseLock( R2511 ),
       //.io_requests_6_7_grant(  )
       .io_requests_6_7_request( T2510 ),
       //.io_requests_6_7_priorityLevel(  )
       .io_requests_6_6_releaseLock( R2506 ),
       //.io_requests_6_6_grant(  )
       .io_requests_6_6_request( T2505 ),
       //.io_requests_6_6_priorityLevel(  )
       .io_requests_6_5_releaseLock( R2501 ),
       //.io_requests_6_5_grant(  )
       .io_requests_6_5_request( T2500 ),
       //.io_requests_6_5_priorityLevel(  )
       .io_requests_6_4_releaseLock( R2496 ),
       //.io_requests_6_4_grant(  )
       .io_requests_6_4_request( T2495 ),
       //.io_requests_6_4_priorityLevel(  )
       .io_requests_6_3_releaseLock( R2491 ),
       //.io_requests_6_3_grant(  )
       .io_requests_6_3_request( T2490 ),
       //.io_requests_6_3_priorityLevel(  )
       .io_requests_6_2_releaseLock( R2486 ),
       //.io_requests_6_2_grant(  )
       .io_requests_6_2_request( T2485 ),
       //.io_requests_6_2_priorityLevel(  )
       .io_requests_6_1_releaseLock( R2481 ),
       //.io_requests_6_1_grant(  )
       .io_requests_6_1_request( T2480 ),
       //.io_requests_6_1_priorityLevel(  )
       .io_requests_6_0_releaseLock( R2476 ),
       //.io_requests_6_0_grant(  )
       .io_requests_6_0_request( T2475 ),
       //.io_requests_6_0_priorityLevel(  )
       .io_requests_5_9_releaseLock( R2471 ),
       //.io_requests_5_9_grant(  )
       .io_requests_5_9_request( T2470 ),
       //.io_requests_5_9_priorityLevel(  )
       .io_requests_5_8_releaseLock( R2466 ),
       //.io_requests_5_8_grant(  )
       .io_requests_5_8_request( T2465 ),
       //.io_requests_5_8_priorityLevel(  )
       .io_requests_5_7_releaseLock( R2461 ),
       //.io_requests_5_7_grant(  )
       .io_requests_5_7_request( T2460 ),
       //.io_requests_5_7_priorityLevel(  )
       .io_requests_5_6_releaseLock( R2456 ),
       //.io_requests_5_6_grant(  )
       .io_requests_5_6_request( T2455 ),
       //.io_requests_5_6_priorityLevel(  )
       .io_requests_5_5_releaseLock( R2451 ),
       //.io_requests_5_5_grant(  )
       .io_requests_5_5_request( T2450 ),
       //.io_requests_5_5_priorityLevel(  )
       .io_requests_5_4_releaseLock( R2446 ),
       //.io_requests_5_4_grant(  )
       .io_requests_5_4_request( T2445 ),
       //.io_requests_5_4_priorityLevel(  )
       .io_requests_5_3_releaseLock( R2441 ),
       //.io_requests_5_3_grant(  )
       .io_requests_5_3_request( T2440 ),
       //.io_requests_5_3_priorityLevel(  )
       .io_requests_5_2_releaseLock( R2436 ),
       //.io_requests_5_2_grant(  )
       .io_requests_5_2_request( T2435 ),
       //.io_requests_5_2_priorityLevel(  )
       .io_requests_5_1_releaseLock( R2431 ),
       //.io_requests_5_1_grant(  )
       .io_requests_5_1_request( T2430 ),
       //.io_requests_5_1_priorityLevel(  )
       .io_requests_5_0_releaseLock( R2426 ),
       //.io_requests_5_0_grant(  )
       .io_requests_5_0_request( T2425 ),
       //.io_requests_5_0_priorityLevel(  )
       .io_requests_4_9_releaseLock( R2421 ),
       //.io_requests_4_9_grant(  )
       .io_requests_4_9_request( T2420 ),
       //.io_requests_4_9_priorityLevel(  )
       .io_requests_4_8_releaseLock( R2416 ),
       //.io_requests_4_8_grant(  )
       .io_requests_4_8_request( T2415 ),
       //.io_requests_4_8_priorityLevel(  )
       .io_requests_4_7_releaseLock( R2411 ),
       //.io_requests_4_7_grant(  )
       .io_requests_4_7_request( T2410 ),
       //.io_requests_4_7_priorityLevel(  )
       .io_requests_4_6_releaseLock( R2406 ),
       //.io_requests_4_6_grant(  )
       .io_requests_4_6_request( T2405 ),
       //.io_requests_4_6_priorityLevel(  )
       .io_requests_4_5_releaseLock( R2401 ),
       //.io_requests_4_5_grant(  )
       .io_requests_4_5_request( T2400 ),
       //.io_requests_4_5_priorityLevel(  )
       .io_requests_4_4_releaseLock( R2396 ),
       //.io_requests_4_4_grant(  )
       .io_requests_4_4_request( T2395 ),
       //.io_requests_4_4_priorityLevel(  )
       .io_requests_4_3_releaseLock( R2391 ),
       //.io_requests_4_3_grant(  )
       .io_requests_4_3_request( T2390 ),
       //.io_requests_4_3_priorityLevel(  )
       .io_requests_4_2_releaseLock( R2386 ),
       //.io_requests_4_2_grant(  )
       .io_requests_4_2_request( T2385 ),
       //.io_requests_4_2_priorityLevel(  )
       .io_requests_4_1_releaseLock( R2381 ),
       //.io_requests_4_1_grant(  )
       .io_requests_4_1_request( T2380 ),
       //.io_requests_4_1_priorityLevel(  )
       .io_requests_4_0_releaseLock( R2376 ),
       //.io_requests_4_0_grant(  )
       .io_requests_4_0_request( T2375 ),
       //.io_requests_4_0_priorityLevel(  )
       .io_requests_3_9_releaseLock( R2371 ),
       //.io_requests_3_9_grant(  )
       .io_requests_3_9_request( T2370 ),
       //.io_requests_3_9_priorityLevel(  )
       .io_requests_3_8_releaseLock( R2366 ),
       //.io_requests_3_8_grant(  )
       .io_requests_3_8_request( T2365 ),
       //.io_requests_3_8_priorityLevel(  )
       .io_requests_3_7_releaseLock( R2361 ),
       //.io_requests_3_7_grant(  )
       .io_requests_3_7_request( T2360 ),
       //.io_requests_3_7_priorityLevel(  )
       .io_requests_3_6_releaseLock( R2356 ),
       //.io_requests_3_6_grant(  )
       .io_requests_3_6_request( T2355 ),
       //.io_requests_3_6_priorityLevel(  )
       .io_requests_3_5_releaseLock( R2351 ),
       //.io_requests_3_5_grant(  )
       .io_requests_3_5_request( T2350 ),
       //.io_requests_3_5_priorityLevel(  )
       .io_requests_3_4_releaseLock( R2346 ),
       //.io_requests_3_4_grant(  )
       .io_requests_3_4_request( T2345 ),
       //.io_requests_3_4_priorityLevel(  )
       .io_requests_3_3_releaseLock( R2341 ),
       //.io_requests_3_3_grant(  )
       .io_requests_3_3_request( T2340 ),
       //.io_requests_3_3_priorityLevel(  )
       .io_requests_3_2_releaseLock( R2336 ),
       //.io_requests_3_2_grant(  )
       .io_requests_3_2_request( T2335 ),
       //.io_requests_3_2_priorityLevel(  )
       .io_requests_3_1_releaseLock( R2331 ),
       //.io_requests_3_1_grant(  )
       .io_requests_3_1_request( T2330 ),
       //.io_requests_3_1_priorityLevel(  )
       .io_requests_3_0_releaseLock( R2326 ),
       //.io_requests_3_0_grant(  )
       .io_requests_3_0_request( T2325 ),
       //.io_requests_3_0_priorityLevel(  )
       .io_requests_2_9_releaseLock( R2321 ),
       //.io_requests_2_9_grant(  )
       .io_requests_2_9_request( T2320 ),
       //.io_requests_2_9_priorityLevel(  )
       .io_requests_2_8_releaseLock( R2316 ),
       //.io_requests_2_8_grant(  )
       .io_requests_2_8_request( T2315 ),
       //.io_requests_2_8_priorityLevel(  )
       .io_requests_2_7_releaseLock( R2311 ),
       //.io_requests_2_7_grant(  )
       .io_requests_2_7_request( T2310 ),
       //.io_requests_2_7_priorityLevel(  )
       .io_requests_2_6_releaseLock( R2306 ),
       //.io_requests_2_6_grant(  )
       .io_requests_2_6_request( T2305 ),
       //.io_requests_2_6_priorityLevel(  )
       .io_requests_2_5_releaseLock( R2301 ),
       //.io_requests_2_5_grant(  )
       .io_requests_2_5_request( T2300 ),
       //.io_requests_2_5_priorityLevel(  )
       .io_requests_2_4_releaseLock( R2296 ),
       //.io_requests_2_4_grant(  )
       .io_requests_2_4_request( T2295 ),
       //.io_requests_2_4_priorityLevel(  )
       .io_requests_2_3_releaseLock( R2291 ),
       //.io_requests_2_3_grant(  )
       .io_requests_2_3_request( T2290 ),
       //.io_requests_2_3_priorityLevel(  )
       .io_requests_2_2_releaseLock( R2286 ),
       //.io_requests_2_2_grant(  )
       .io_requests_2_2_request( T2285 ),
       //.io_requests_2_2_priorityLevel(  )
       .io_requests_2_1_releaseLock( R2281 ),
       //.io_requests_2_1_grant(  )
       .io_requests_2_1_request( T2280 ),
       //.io_requests_2_1_priorityLevel(  )
       .io_requests_2_0_releaseLock( R2276 ),
       //.io_requests_2_0_grant(  )
       .io_requests_2_0_request( T2275 ),
       //.io_requests_2_0_priorityLevel(  )
       .io_requests_1_9_releaseLock( R2271 ),
       //.io_requests_1_9_grant(  )
       .io_requests_1_9_request( T2270 ),
       //.io_requests_1_9_priorityLevel(  )
       .io_requests_1_8_releaseLock( R2266 ),
       //.io_requests_1_8_grant(  )
       .io_requests_1_8_request( T2265 ),
       //.io_requests_1_8_priorityLevel(  )
       .io_requests_1_7_releaseLock( R2261 ),
       //.io_requests_1_7_grant(  )
       .io_requests_1_7_request( T2260 ),
       //.io_requests_1_7_priorityLevel(  )
       .io_requests_1_6_releaseLock( R2256 ),
       //.io_requests_1_6_grant(  )
       .io_requests_1_6_request( T2255 ),
       //.io_requests_1_6_priorityLevel(  )
       .io_requests_1_5_releaseLock( R2251 ),
       //.io_requests_1_5_grant(  )
       .io_requests_1_5_request( T2250 ),
       //.io_requests_1_5_priorityLevel(  )
       .io_requests_1_4_releaseLock( R2246 ),
       //.io_requests_1_4_grant(  )
       .io_requests_1_4_request( T2245 ),
       //.io_requests_1_4_priorityLevel(  )
       .io_requests_1_3_releaseLock( R2241 ),
       //.io_requests_1_3_grant(  )
       .io_requests_1_3_request( T2240 ),
       //.io_requests_1_3_priorityLevel(  )
       .io_requests_1_2_releaseLock( R2236 ),
       //.io_requests_1_2_grant(  )
       .io_requests_1_2_request( T2235 ),
       //.io_requests_1_2_priorityLevel(  )
       .io_requests_1_1_releaseLock( R2231 ),
       //.io_requests_1_1_grant(  )
       .io_requests_1_1_request( T2230 ),
       //.io_requests_1_1_priorityLevel(  )
       .io_requests_1_0_releaseLock( R2226 ),
       //.io_requests_1_0_grant(  )
       .io_requests_1_0_request( T2225 ),
       //.io_requests_1_0_priorityLevel(  )
       .io_requests_0_9_releaseLock( R2221 ),
       //.io_requests_0_9_grant(  )
       .io_requests_0_9_request( T2220 ),
       //.io_requests_0_9_priorityLevel(  )
       .io_requests_0_8_releaseLock( R2216 ),
       //.io_requests_0_8_grant(  )
       .io_requests_0_8_request( T2215 ),
       //.io_requests_0_8_priorityLevel(  )
       .io_requests_0_7_releaseLock( R2211 ),
       //.io_requests_0_7_grant(  )
       .io_requests_0_7_request( T2210 ),
       //.io_requests_0_7_priorityLevel(  )
       .io_requests_0_6_releaseLock( R2206 ),
       //.io_requests_0_6_grant(  )
       .io_requests_0_6_request( T2205 ),
       //.io_requests_0_6_priorityLevel(  )
       .io_requests_0_5_releaseLock( R2201 ),
       //.io_requests_0_5_grant(  )
       .io_requests_0_5_request( T2200 ),
       //.io_requests_0_5_priorityLevel(  )
       .io_requests_0_4_releaseLock( R2196 ),
       //.io_requests_0_4_grant(  )
       .io_requests_0_4_request( T2195 ),
       //.io_requests_0_4_priorityLevel(  )
       .io_requests_0_3_releaseLock( R2191 ),
       //.io_requests_0_3_grant(  )
       .io_requests_0_3_request( T2190 ),
       //.io_requests_0_3_priorityLevel(  )
       .io_requests_0_2_releaseLock( R2186 ),
       //.io_requests_0_2_grant(  )
       .io_requests_0_2_request( T2185 ),
       //.io_requests_0_2_priorityLevel(  )
       .io_requests_0_1_releaseLock( R2181 ),
       //.io_requests_0_1_grant(  )
       .io_requests_0_1_request( T2180 ),
       //.io_requests_0_1_priorityLevel(  )
       .io_requests_0_0_releaseLock( R2176 ),
       //.io_requests_0_0_grant(  )
       .io_requests_0_0_request( T2175 ),
       //.io_requests_0_0_priorityLevel(  )
       .io_resources_9_ready( T2173 ),
       .io_resources_9_valid( vcAllocator_io_resources_9_valid ),
       .io_resources_8_ready( T2171 ),
       .io_resources_8_valid( vcAllocator_io_resources_8_valid ),
       .io_resources_7_ready( T2169 ),
       .io_resources_7_valid( vcAllocator_io_resources_7_valid ),
       .io_resources_6_ready( T2167 ),
       .io_resources_6_valid( vcAllocator_io_resources_6_valid ),
       .io_resources_5_ready( T2165 ),
       .io_resources_5_valid( vcAllocator_io_resources_5_valid ),
       .io_resources_4_ready( T2163 ),
       .io_resources_4_valid( vcAllocator_io_resources_4_valid ),
       .io_resources_3_ready( T2161 ),
       .io_resources_3_valid( vcAllocator_io_resources_3_valid ),
       .io_resources_2_ready( T2159 ),
       .io_resources_2_valid( vcAllocator_io_resources_2_valid ),
       .io_resources_1_ready( T2157 ),
       .io_resources_1_valid( vcAllocator_io_resources_1_valid ),
       .io_resources_0_ready( T2155 ),
       .io_resources_0_valid( vcAllocator_io_resources_0_valid ),
       .io_chosens_9( vcAllocator_io_chosens_9 ),
       .io_chosens_8( vcAllocator_io_chosens_8 ),
       .io_chosens_7( vcAllocator_io_chosens_7 ),
       .io_chosens_6( vcAllocator_io_chosens_6 ),
       .io_chosens_5( vcAllocator_io_chosens_5 ),
       .io_chosens_4( vcAllocator_io_chosens_4 ),
       .io_chosens_3( vcAllocator_io_chosens_3 ),
       .io_chosens_2( vcAllocator_io_chosens_2 ),
       .io_chosens_1( vcAllocator_io_chosens_1 ),
       .io_chosens_0( vcAllocator_io_chosens_0 )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign vcAllocator.io_requests_9_9_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_9_8_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_9_7_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_9_6_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_9_5_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_9_4_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_9_3_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_9_2_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_9_1_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_9_0_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_8_9_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_8_8_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_8_7_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_8_6_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_8_5_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_8_4_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_8_3_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_8_2_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_8_1_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_8_0_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_7_9_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_7_8_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_7_7_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_7_6_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_7_5_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_7_4_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_7_3_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_7_2_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_7_1_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_7_0_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_6_9_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_6_8_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_6_7_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_6_6_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_6_5_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_6_4_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_6_3_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_6_2_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_6_1_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_6_0_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_5_9_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_5_8_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_5_7_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_5_6_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_5_5_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_5_4_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_5_3_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_5_2_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_5_1_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_5_0_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_4_9_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_4_8_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_4_7_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_4_6_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_4_5_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_4_4_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_4_3_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_4_2_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_4_1_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_4_0_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_3_9_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_3_8_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_3_7_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_3_6_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_3_5_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_3_4_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_3_3_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_3_2_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_3_1_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_3_0_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_2_9_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_2_8_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_2_7_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_2_6_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_2_5_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_2_4_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_2_3_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_2_2_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_2_1_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_2_0_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_1_9_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_1_8_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_1_7_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_1_6_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_1_5_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_1_4_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_1_3_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_1_2_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_1_1_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_1_0_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_0_9_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_0_8_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_0_7_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_0_6_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_0_5_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_0_4_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_0_3_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_0_2_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_0_1_priorityLevel = {1{1'b0}};
    assign vcAllocator.io_requests_0_0_priorityLevel = {1{1'b0}};
// synthesis translate_on
`endif
  VCRouterOutputStateManagement VCRouterOutputStateManagement(.clk(clk), .reset(reset),
       .io_swAllocGranted( T2094 ),
       .io_creditsAvail( T2092 ),
       .io_currentState( VCRouterOutputStateManagement_io_currentState )
  );
  VCRouterOutputStateManagement VCRouterOutputStateManagement_1(.clk(clk), .reset(reset),
       .io_swAllocGranted( T2031 ),
       .io_creditsAvail( T2029 ),
       .io_currentState( VCRouterOutputStateManagement_1_io_currentState )
  );
  VCRouterOutputStateManagement VCRouterOutputStateManagement_2(.clk(clk), .reset(reset),
       .io_swAllocGranted( T1968 ),
       .io_creditsAvail( T1966 ),
       .io_currentState( VCRouterOutputStateManagement_2_io_currentState )
  );
  VCRouterOutputStateManagement VCRouterOutputStateManagement_3(.clk(clk), .reset(reset),
       .io_swAllocGranted( T1905 ),
       .io_creditsAvail( T1903 ),
       .io_currentState( VCRouterOutputStateManagement_3_io_currentState )
  );
  VCRouterOutputStateManagement VCRouterOutputStateManagement_4(.clk(clk), .reset(reset),
       .io_swAllocGranted( T1722 ),
       .io_creditsAvail( T1720 ),
       .io_currentState( VCRouterOutputStateManagement_4_io_currentState )
  );
  CreditGen CreditGen(
       .io_outCredit_grant( CreditGen_io_outCredit_grant ),
       .io_inGrant( T1710 )
  );
  RouterRegFile RouterRegFile(.clk(clk), .reset(reset),
       .io_writeData( T1708 ),
       .io_writeEnable( T1705 ),
       //.io_full(  )
       .io_readData( RouterRegFile_io_readData ),
       .io_readValid( RouterRegFile_io_readValid ),
       .io_readIncrement( T1692 ),
       .io_writePipelineReg_2( RouterRegFile_io_readPipelineReg_1 ),
       .io_writePipelineReg_1( RouterRegFile_io_readPipelineReg_0 ),
       .io_writePipelineReg_0( T3181 ),
       .io_wePipelineReg_2( T1681 ),
       .io_wePipelineReg_1( T1678 ),
       .io_wePipelineReg_0( T1676 ),
       //.io_readPipelineReg_2(  )
       .io_readPipelineReg_1( RouterRegFile_io_readPipelineReg_1 ),
       .io_readPipelineReg_0( RouterRegFile_io_readPipelineReg_0 ),
       //.io_rvPipelineReg_2(  )
       .io_rvPipelineReg_1( RouterRegFile_io_rvPipelineReg_1 ),
       .io_rvPipelineReg_0( RouterRegFile_io_rvPipelineReg_0 )
  );
  RouterBuffer RouterBuffer(.clk(clk), .reset(reset),
       .io_enq_ready( RouterBuffer_io_enq_ready ),
       .io_enq_valid( T1675 ),
       .io_enq_bits_x( io_inChannels_0_flit_x ),
       .io_deq_ready( T1656 ),
       .io_deq_valid( RouterBuffer_io_deq_valid ),
       .io_deq_bits_x( RouterBuffer_io_deq_bits_x )
  );
  CMeshDOR_2 CMeshDOR(
       .io_inHeadFlit_packetID( T1655 ),
       .io_inHeadFlit_isTail( T1654 ),
       .io_inHeadFlit_vcPort( T1653 ),
       .io_inHeadFlit_packetType( T1652 ),
       .io_inHeadFlit_destination_2( T1651 ),
       .io_inHeadFlit_destination_1( T1650 ),
       .io_inHeadFlit_destination_0( T1649 ),
       .io_inHeadFlit_priorityLevel( T1646 ),
       .io_outHeadFlit_packetID( CMeshDOR_io_outHeadFlit_packetID ),
       .io_outHeadFlit_isTail( CMeshDOR_io_outHeadFlit_isTail ),
       .io_outHeadFlit_vcPort( CMeshDOR_io_outHeadFlit_vcPort ),
       .io_outHeadFlit_packetType( CMeshDOR_io_outHeadFlit_packetType ),
       .io_outHeadFlit_destination_2( CMeshDOR_io_outHeadFlit_destination_2 ),
       .io_outHeadFlit_destination_1( CMeshDOR_io_outHeadFlit_destination_1 ),
       .io_outHeadFlit_destination_0( CMeshDOR_io_outHeadFlit_destination_0 ),
       .io_outHeadFlit_priorityLevel( CMeshDOR_io_outHeadFlit_priorityLevel ),
       .io_result( CMeshDOR_io_result ),
       .io_vcsAvailable_4( CMeshDOR_io_vcsAvailable_4 ),
       .io_vcsAvailable_3( CMeshDOR_io_vcsAvailable_3 ),
       .io_vcsAvailable_2( CMeshDOR_io_vcsAvailable_2 ),
       .io_vcsAvailable_1( CMeshDOR_io_vcsAvailable_1 ),
       .io_vcsAvailable_0( CMeshDOR_io_vcsAvailable_0 )
  );
  VCRouterStateManagement VCRouterStateManagement(.clk(clk), .reset(reset),
       .io_inputBufferValid( RouterBuffer_io_deq_valid ),
       .io_routingComplete( R1645 ),
       .io_inputBufferIsTail( T1636 ),
       .io_vcAllocGranted( vcAllocator_io_resources_0_valid ),
       .io_swAllocGranted( T1616 ),
       .io_creditsAvail( T1597 ),
       .io_outputReady( T1584 ),
       .io_currentState( VCRouterStateManagement_io_currentState )
  );
  ReplaceVCPort ReplaceVCPort(
       .io_oldFlit_x( T1582 ),
       .io_newVCPort( T3175 ),
       .io_newFlit_x( ReplaceVCPort_io_newFlit_x )
  );
  Flit2FlitBundle Flit2FlitBundle(
       .io_inFlit_x( T1576 )
       //.io_outHead_packetID(  )
       //.io_outHead_isTail(  )
       //.io_outHead_vcPort(  )
       //.io_outHead_packetType(  )
       //.io_outHead_destination_2(  )
       //.io_outHead_destination_1(  )
       //.io_outHead_destination_0(  )
       //.io_outHead_priorityLevel(  )
       //.io_outBody_packetID(  )
       //.io_outBody_isTail(  )
       //.io_outBody_vcPort(  )
       //.io_outBody_flitID(  )
       //.io_outBody_payload(  )
  );
  CreditGen CreditGen_1(
       .io_outCredit_grant( CreditGen_1_io_outCredit_grant ),
       .io_inGrant( T1566 )
  );
  RouterRegFile RouterRegFile_1(.clk(clk), .reset(reset),
       .io_writeData( T1564 ),
       .io_writeEnable( T1561 ),
       //.io_full(  )
       .io_readData( RouterRegFile_1_io_readData ),
       .io_readValid( RouterRegFile_1_io_readValid ),
       .io_readIncrement( T1548 ),
       .io_writePipelineReg_2( RouterRegFile_1_io_readPipelineReg_1 ),
       .io_writePipelineReg_1( RouterRegFile_1_io_readPipelineReg_0 ),
       .io_writePipelineReg_0( T3174 ),
       .io_wePipelineReg_2( T1537 ),
       .io_wePipelineReg_1( T1534 ),
       .io_wePipelineReg_0( T1532 ),
       //.io_readPipelineReg_2(  )
       .io_readPipelineReg_1( RouterRegFile_1_io_readPipelineReg_1 ),
       .io_readPipelineReg_0( RouterRegFile_1_io_readPipelineReg_0 ),
       //.io_rvPipelineReg_2(  )
       .io_rvPipelineReg_1( RouterRegFile_1_io_rvPipelineReg_1 ),
       .io_rvPipelineReg_0( RouterRegFile_1_io_rvPipelineReg_0 )
  );
  RouterBuffer RouterBuffer_1(.clk(clk), .reset(reset),
       .io_enq_ready( RouterBuffer_1_io_enq_ready ),
       .io_enq_valid( T1531 ),
       .io_enq_bits_x( io_inChannels_0_flit_x ),
       .io_deq_ready( T1512 ),
       .io_deq_valid( RouterBuffer_1_io_deq_valid ),
       .io_deq_bits_x( RouterBuffer_1_io_deq_bits_x )
  );
  CMeshDOR_2 CMeshDOR_1(
       .io_inHeadFlit_packetID( T1511 ),
       .io_inHeadFlit_isTail( T1510 ),
       .io_inHeadFlit_vcPort( T1509 ),
       .io_inHeadFlit_packetType( T1508 ),
       .io_inHeadFlit_destination_2( T1507 ),
       .io_inHeadFlit_destination_1( T1506 ),
       .io_inHeadFlit_destination_0( T1505 ),
       .io_inHeadFlit_priorityLevel( T1502 ),
       .io_outHeadFlit_packetID( CMeshDOR_1_io_outHeadFlit_packetID ),
       .io_outHeadFlit_isTail( CMeshDOR_1_io_outHeadFlit_isTail ),
       .io_outHeadFlit_vcPort( CMeshDOR_1_io_outHeadFlit_vcPort ),
       .io_outHeadFlit_packetType( CMeshDOR_1_io_outHeadFlit_packetType ),
       .io_outHeadFlit_destination_2( CMeshDOR_1_io_outHeadFlit_destination_2 ),
       .io_outHeadFlit_destination_1( CMeshDOR_1_io_outHeadFlit_destination_1 ),
       .io_outHeadFlit_destination_0( CMeshDOR_1_io_outHeadFlit_destination_0 ),
       .io_outHeadFlit_priorityLevel( CMeshDOR_1_io_outHeadFlit_priorityLevel ),
       .io_result( CMeshDOR_1_io_result ),
       .io_vcsAvailable_4( CMeshDOR_1_io_vcsAvailable_4 ),
       .io_vcsAvailable_3( CMeshDOR_1_io_vcsAvailable_3 ),
       .io_vcsAvailable_2( CMeshDOR_1_io_vcsAvailable_2 ),
       .io_vcsAvailable_1( CMeshDOR_1_io_vcsAvailable_1 ),
       .io_vcsAvailable_0( CMeshDOR_1_io_vcsAvailable_0 )
  );
  VCRouterStateManagement VCRouterStateManagement_1(.clk(clk), .reset(reset),
       .io_inputBufferValid( RouterBuffer_1_io_deq_valid ),
       .io_routingComplete( R1501 ),
       .io_inputBufferIsTail( T1492 ),
       .io_vcAllocGranted( vcAllocator_io_resources_1_valid ),
       .io_swAllocGranted( T1472 ),
       .io_creditsAvail( T1453 ),
       .io_outputReady( T1440 ),
       .io_currentState( VCRouterStateManagement_1_io_currentState )
  );
  ReplaceVCPort ReplaceVCPort_1(
       .io_oldFlit_x( T1438 ),
       .io_newVCPort( T3168 ),
       .io_newFlit_x( ReplaceVCPort_1_io_newFlit_x )
  );
  Flit2FlitBundle Flit2FlitBundle_1(
       .io_inFlit_x( T1432 )
       //.io_outHead_packetID(  )
       //.io_outHead_isTail(  )
       //.io_outHead_vcPort(  )
       //.io_outHead_packetType(  )
       //.io_outHead_destination_2(  )
       //.io_outHead_destination_1(  )
       //.io_outHead_destination_0(  )
       //.io_outHead_priorityLevel(  )
       //.io_outBody_packetID(  )
       //.io_outBody_isTail(  )
       //.io_outBody_vcPort(  )
       //.io_outBody_flitID(  )
       //.io_outBody_payload(  )
  );
  CreditGen CreditGen_2(
       .io_outCredit_grant( CreditGen_2_io_outCredit_grant ),
       .io_inGrant( T1422 )
  );
  RouterRegFile RouterRegFile_2(.clk(clk), .reset(reset),
       .io_writeData( T1420 ),
       .io_writeEnable( T1417 ),
       //.io_full(  )
       .io_readData( RouterRegFile_2_io_readData ),
       .io_readValid( RouterRegFile_2_io_readValid ),
       .io_readIncrement( T1404 ),
       .io_writePipelineReg_2( RouterRegFile_2_io_readPipelineReg_1 ),
       .io_writePipelineReg_1( RouterRegFile_2_io_readPipelineReg_0 ),
       .io_writePipelineReg_0( T3167 ),
       .io_wePipelineReg_2( T1393 ),
       .io_wePipelineReg_1( T1390 ),
       .io_wePipelineReg_0( T1388 ),
       //.io_readPipelineReg_2(  )
       .io_readPipelineReg_1( RouterRegFile_2_io_readPipelineReg_1 ),
       .io_readPipelineReg_0( RouterRegFile_2_io_readPipelineReg_0 ),
       //.io_rvPipelineReg_2(  )
       .io_rvPipelineReg_1( RouterRegFile_2_io_rvPipelineReg_1 ),
       .io_rvPipelineReg_0( RouterRegFile_2_io_rvPipelineReg_0 )
  );
  RouterBuffer RouterBuffer_2(.clk(clk), .reset(reset),
       .io_enq_ready( RouterBuffer_2_io_enq_ready ),
       .io_enq_valid( T1387 ),
       .io_enq_bits_x( io_inChannels_1_flit_x ),
       .io_deq_ready( T1368 ),
       .io_deq_valid( RouterBuffer_2_io_deq_valid ),
       .io_deq_bits_x( RouterBuffer_2_io_deq_bits_x )
  );
  CMeshDOR_2 CMeshDOR_2(
       .io_inHeadFlit_packetID( T1367 ),
       .io_inHeadFlit_isTail( T1366 ),
       .io_inHeadFlit_vcPort( T1365 ),
       .io_inHeadFlit_packetType( T1364 ),
       .io_inHeadFlit_destination_2( T1363 ),
       .io_inHeadFlit_destination_1( T1362 ),
       .io_inHeadFlit_destination_0( T1361 ),
       .io_inHeadFlit_priorityLevel( T1358 ),
       .io_outHeadFlit_packetID( CMeshDOR_2_io_outHeadFlit_packetID ),
       .io_outHeadFlit_isTail( CMeshDOR_2_io_outHeadFlit_isTail ),
       .io_outHeadFlit_vcPort( CMeshDOR_2_io_outHeadFlit_vcPort ),
       .io_outHeadFlit_packetType( CMeshDOR_2_io_outHeadFlit_packetType ),
       .io_outHeadFlit_destination_2( CMeshDOR_2_io_outHeadFlit_destination_2 ),
       .io_outHeadFlit_destination_1( CMeshDOR_2_io_outHeadFlit_destination_1 ),
       .io_outHeadFlit_destination_0( CMeshDOR_2_io_outHeadFlit_destination_0 ),
       .io_outHeadFlit_priorityLevel( CMeshDOR_2_io_outHeadFlit_priorityLevel ),
       .io_result( CMeshDOR_2_io_result ),
       .io_vcsAvailable_4( CMeshDOR_2_io_vcsAvailable_4 ),
       .io_vcsAvailable_3( CMeshDOR_2_io_vcsAvailable_3 ),
       .io_vcsAvailable_2( CMeshDOR_2_io_vcsAvailable_2 ),
       .io_vcsAvailable_1( CMeshDOR_2_io_vcsAvailable_1 ),
       .io_vcsAvailable_0( CMeshDOR_2_io_vcsAvailable_0 )
  );
  VCRouterStateManagement VCRouterStateManagement_2(.clk(clk), .reset(reset),
       .io_inputBufferValid( RouterBuffer_2_io_deq_valid ),
       .io_routingComplete( R1357 ),
       .io_inputBufferIsTail( T1348 ),
       .io_vcAllocGranted( vcAllocator_io_resources_2_valid ),
       .io_swAllocGranted( T1328 ),
       .io_creditsAvail( T1309 ),
       .io_outputReady( T1296 ),
       .io_currentState( VCRouterStateManagement_2_io_currentState )
  );
  ReplaceVCPort ReplaceVCPort_2(
       .io_oldFlit_x( T1294 ),
       .io_newVCPort( T3161 ),
       .io_newFlit_x( ReplaceVCPort_2_io_newFlit_x )
  );
  Flit2FlitBundle Flit2FlitBundle_2(
       .io_inFlit_x( T1288 )
       //.io_outHead_packetID(  )
       //.io_outHead_isTail(  )
       //.io_outHead_vcPort(  )
       //.io_outHead_packetType(  )
       //.io_outHead_destination_2(  )
       //.io_outHead_destination_1(  )
       //.io_outHead_destination_0(  )
       //.io_outHead_priorityLevel(  )
       //.io_outBody_packetID(  )
       //.io_outBody_isTail(  )
       //.io_outBody_vcPort(  )
       //.io_outBody_flitID(  )
       //.io_outBody_payload(  )
  );
  CreditGen CreditGen_3(
       .io_outCredit_grant( CreditGen_3_io_outCredit_grant ),
       .io_inGrant( T1278 )
  );
  RouterRegFile RouterRegFile_3(.clk(clk), .reset(reset),
       .io_writeData( T1276 ),
       .io_writeEnable( T1273 ),
       //.io_full(  )
       .io_readData( RouterRegFile_3_io_readData ),
       .io_readValid( RouterRegFile_3_io_readValid ),
       .io_readIncrement( T1260 ),
       .io_writePipelineReg_2( RouterRegFile_3_io_readPipelineReg_1 ),
       .io_writePipelineReg_1( RouterRegFile_3_io_readPipelineReg_0 ),
       .io_writePipelineReg_0( T3160 ),
       .io_wePipelineReg_2( T1249 ),
       .io_wePipelineReg_1( T1246 ),
       .io_wePipelineReg_0( T1244 ),
       //.io_readPipelineReg_2(  )
       .io_readPipelineReg_1( RouterRegFile_3_io_readPipelineReg_1 ),
       .io_readPipelineReg_0( RouterRegFile_3_io_readPipelineReg_0 ),
       //.io_rvPipelineReg_2(  )
       .io_rvPipelineReg_1( RouterRegFile_3_io_rvPipelineReg_1 ),
       .io_rvPipelineReg_0( RouterRegFile_3_io_rvPipelineReg_0 )
  );
  RouterBuffer RouterBuffer_3(.clk(clk), .reset(reset),
       .io_enq_ready( RouterBuffer_3_io_enq_ready ),
       .io_enq_valid( T1243 ),
       .io_enq_bits_x( io_inChannels_1_flit_x ),
       .io_deq_ready( T1224 ),
       .io_deq_valid( RouterBuffer_3_io_deq_valid ),
       .io_deq_bits_x( RouterBuffer_3_io_deq_bits_x )
  );
  CMeshDOR_2 CMeshDOR_3(
       .io_inHeadFlit_packetID( T1223 ),
       .io_inHeadFlit_isTail( T1222 ),
       .io_inHeadFlit_vcPort( T1221 ),
       .io_inHeadFlit_packetType( T1220 ),
       .io_inHeadFlit_destination_2( T1219 ),
       .io_inHeadFlit_destination_1( T1218 ),
       .io_inHeadFlit_destination_0( T1217 ),
       .io_inHeadFlit_priorityLevel( T1214 ),
       .io_outHeadFlit_packetID( CMeshDOR_3_io_outHeadFlit_packetID ),
       .io_outHeadFlit_isTail( CMeshDOR_3_io_outHeadFlit_isTail ),
       .io_outHeadFlit_vcPort( CMeshDOR_3_io_outHeadFlit_vcPort ),
       .io_outHeadFlit_packetType( CMeshDOR_3_io_outHeadFlit_packetType ),
       .io_outHeadFlit_destination_2( CMeshDOR_3_io_outHeadFlit_destination_2 ),
       .io_outHeadFlit_destination_1( CMeshDOR_3_io_outHeadFlit_destination_1 ),
       .io_outHeadFlit_destination_0( CMeshDOR_3_io_outHeadFlit_destination_0 ),
       .io_outHeadFlit_priorityLevel( CMeshDOR_3_io_outHeadFlit_priorityLevel ),
       .io_result( CMeshDOR_3_io_result ),
       .io_vcsAvailable_4( CMeshDOR_3_io_vcsAvailable_4 ),
       .io_vcsAvailable_3( CMeshDOR_3_io_vcsAvailable_3 ),
       .io_vcsAvailable_2( CMeshDOR_3_io_vcsAvailable_2 ),
       .io_vcsAvailable_1( CMeshDOR_3_io_vcsAvailable_1 ),
       .io_vcsAvailable_0( CMeshDOR_3_io_vcsAvailable_0 )
  );
  VCRouterStateManagement VCRouterStateManagement_3(.clk(clk), .reset(reset),
       .io_inputBufferValid( RouterBuffer_3_io_deq_valid ),
       .io_routingComplete( R1213 ),
       .io_inputBufferIsTail( T1204 ),
       .io_vcAllocGranted( vcAllocator_io_resources_3_valid ),
       .io_swAllocGranted( T1184 ),
       .io_creditsAvail( T1165 ),
       .io_outputReady( T1152 ),
       .io_currentState( VCRouterStateManagement_3_io_currentState )
  );
  ReplaceVCPort ReplaceVCPort_3(
       .io_oldFlit_x( T1150 ),
       .io_newVCPort( T3154 ),
       .io_newFlit_x( ReplaceVCPort_3_io_newFlit_x )
  );
  Flit2FlitBundle Flit2FlitBundle_3(
       .io_inFlit_x( T1144 )
       //.io_outHead_packetID(  )
       //.io_outHead_isTail(  )
       //.io_outHead_vcPort(  )
       //.io_outHead_packetType(  )
       //.io_outHead_destination_2(  )
       //.io_outHead_destination_1(  )
       //.io_outHead_destination_0(  )
       //.io_outHead_priorityLevel(  )
       //.io_outBody_packetID(  )
       //.io_outBody_isTail(  )
       //.io_outBody_vcPort(  )
       //.io_outBody_flitID(  )
       //.io_outBody_payload(  )
  );
  CreditGen CreditGen_4(
       .io_outCredit_grant( CreditGen_4_io_outCredit_grant ),
       .io_inGrant( T1134 )
  );
  RouterRegFile RouterRegFile_4(.clk(clk), .reset(reset),
       .io_writeData( T1132 ),
       .io_writeEnable( T1129 ),
       //.io_full(  )
       .io_readData( RouterRegFile_4_io_readData ),
       .io_readValid( RouterRegFile_4_io_readValid ),
       .io_readIncrement( T1116 ),
       .io_writePipelineReg_2( RouterRegFile_4_io_readPipelineReg_1 ),
       .io_writePipelineReg_1( RouterRegFile_4_io_readPipelineReg_0 ),
       .io_writePipelineReg_0( T3153 ),
       .io_wePipelineReg_2( T1105 ),
       .io_wePipelineReg_1( T1102 ),
       .io_wePipelineReg_0( T1100 ),
       //.io_readPipelineReg_2(  )
       .io_readPipelineReg_1( RouterRegFile_4_io_readPipelineReg_1 ),
       .io_readPipelineReg_0( RouterRegFile_4_io_readPipelineReg_0 ),
       //.io_rvPipelineReg_2(  )
       .io_rvPipelineReg_1( RouterRegFile_4_io_rvPipelineReg_1 ),
       .io_rvPipelineReg_0( RouterRegFile_4_io_rvPipelineReg_0 )
  );
  RouterBuffer RouterBuffer_4(.clk(clk), .reset(reset),
       .io_enq_ready( RouterBuffer_4_io_enq_ready ),
       .io_enq_valid( T1099 ),
       .io_enq_bits_x( io_inChannels_2_flit_x ),
       .io_deq_ready( T1080 ),
       .io_deq_valid( RouterBuffer_4_io_deq_valid ),
       .io_deq_bits_x( RouterBuffer_4_io_deq_bits_x )
  );
  CMeshDOR_2 CMeshDOR_4(
       .io_inHeadFlit_packetID( T1079 ),
       .io_inHeadFlit_isTail( T1078 ),
       .io_inHeadFlit_vcPort( T1077 ),
       .io_inHeadFlit_packetType( T1076 ),
       .io_inHeadFlit_destination_2( T1075 ),
       .io_inHeadFlit_destination_1( T1074 ),
       .io_inHeadFlit_destination_0( T1073 ),
       .io_inHeadFlit_priorityLevel( T1070 ),
       .io_outHeadFlit_packetID( CMeshDOR_4_io_outHeadFlit_packetID ),
       .io_outHeadFlit_isTail( CMeshDOR_4_io_outHeadFlit_isTail ),
       .io_outHeadFlit_vcPort( CMeshDOR_4_io_outHeadFlit_vcPort ),
       .io_outHeadFlit_packetType( CMeshDOR_4_io_outHeadFlit_packetType ),
       .io_outHeadFlit_destination_2( CMeshDOR_4_io_outHeadFlit_destination_2 ),
       .io_outHeadFlit_destination_1( CMeshDOR_4_io_outHeadFlit_destination_1 ),
       .io_outHeadFlit_destination_0( CMeshDOR_4_io_outHeadFlit_destination_0 ),
       .io_outHeadFlit_priorityLevel( CMeshDOR_4_io_outHeadFlit_priorityLevel ),
       .io_result( CMeshDOR_4_io_result ),
       .io_vcsAvailable_4( CMeshDOR_4_io_vcsAvailable_4 ),
       .io_vcsAvailable_3( CMeshDOR_4_io_vcsAvailable_3 ),
       .io_vcsAvailable_2( CMeshDOR_4_io_vcsAvailable_2 ),
       .io_vcsAvailable_1( CMeshDOR_4_io_vcsAvailable_1 ),
       .io_vcsAvailable_0( CMeshDOR_4_io_vcsAvailable_0 )
  );
  VCRouterStateManagement VCRouterStateManagement_4(.clk(clk), .reset(reset),
       .io_inputBufferValid( RouterBuffer_4_io_deq_valid ),
       .io_routingComplete( R1069 ),
       .io_inputBufferIsTail( T1060 ),
       .io_vcAllocGranted( vcAllocator_io_resources_4_valid ),
       .io_swAllocGranted( T1040 ),
       .io_creditsAvail( T1021 ),
       .io_outputReady( T1008 ),
       .io_currentState( VCRouterStateManagement_4_io_currentState )
  );
  ReplaceVCPort ReplaceVCPort_4(
       .io_oldFlit_x( T1006 ),
       .io_newVCPort( T3147 ),
       .io_newFlit_x( ReplaceVCPort_4_io_newFlit_x )
  );
  Flit2FlitBundle Flit2FlitBundle_4(
       .io_inFlit_x( T1000 )
       //.io_outHead_packetID(  )
       //.io_outHead_isTail(  )
       //.io_outHead_vcPort(  )
       //.io_outHead_packetType(  )
       //.io_outHead_destination_2(  )
       //.io_outHead_destination_1(  )
       //.io_outHead_destination_0(  )
       //.io_outHead_priorityLevel(  )
       //.io_outBody_packetID(  )
       //.io_outBody_isTail(  )
       //.io_outBody_vcPort(  )
       //.io_outBody_flitID(  )
       //.io_outBody_payload(  )
  );
  CreditGen CreditGen_5(
       .io_outCredit_grant( CreditGen_5_io_outCredit_grant ),
       .io_inGrant( T990 )
  );
  RouterRegFile RouterRegFile_5(.clk(clk), .reset(reset),
       .io_writeData( T988 ),
       .io_writeEnable( T985 ),
       //.io_full(  )
       .io_readData( RouterRegFile_5_io_readData ),
       .io_readValid( RouterRegFile_5_io_readValid ),
       .io_readIncrement( T972 ),
       .io_writePipelineReg_2( RouterRegFile_5_io_readPipelineReg_1 ),
       .io_writePipelineReg_1( RouterRegFile_5_io_readPipelineReg_0 ),
       .io_writePipelineReg_0( T3146 ),
       .io_wePipelineReg_2( T961 ),
       .io_wePipelineReg_1( T958 ),
       .io_wePipelineReg_0( T956 ),
       //.io_readPipelineReg_2(  )
       .io_readPipelineReg_1( RouterRegFile_5_io_readPipelineReg_1 ),
       .io_readPipelineReg_0( RouterRegFile_5_io_readPipelineReg_0 ),
       //.io_rvPipelineReg_2(  )
       .io_rvPipelineReg_1( RouterRegFile_5_io_rvPipelineReg_1 ),
       .io_rvPipelineReg_0( RouterRegFile_5_io_rvPipelineReg_0 )
  );
  RouterBuffer RouterBuffer_5(.clk(clk), .reset(reset),
       .io_enq_ready( RouterBuffer_5_io_enq_ready ),
       .io_enq_valid( T955 ),
       .io_enq_bits_x( io_inChannels_2_flit_x ),
       .io_deq_ready( T936 ),
       .io_deq_valid( RouterBuffer_5_io_deq_valid ),
       .io_deq_bits_x( RouterBuffer_5_io_deq_bits_x )
  );
  CMeshDOR_2 CMeshDOR_5(
       .io_inHeadFlit_packetID( T935 ),
       .io_inHeadFlit_isTail( T934 ),
       .io_inHeadFlit_vcPort( T933 ),
       .io_inHeadFlit_packetType( T932 ),
       .io_inHeadFlit_destination_2( T931 ),
       .io_inHeadFlit_destination_1( T930 ),
       .io_inHeadFlit_destination_0( T929 ),
       .io_inHeadFlit_priorityLevel( T926 ),
       .io_outHeadFlit_packetID( CMeshDOR_5_io_outHeadFlit_packetID ),
       .io_outHeadFlit_isTail( CMeshDOR_5_io_outHeadFlit_isTail ),
       .io_outHeadFlit_vcPort( CMeshDOR_5_io_outHeadFlit_vcPort ),
       .io_outHeadFlit_packetType( CMeshDOR_5_io_outHeadFlit_packetType ),
       .io_outHeadFlit_destination_2( CMeshDOR_5_io_outHeadFlit_destination_2 ),
       .io_outHeadFlit_destination_1( CMeshDOR_5_io_outHeadFlit_destination_1 ),
       .io_outHeadFlit_destination_0( CMeshDOR_5_io_outHeadFlit_destination_0 ),
       .io_outHeadFlit_priorityLevel( CMeshDOR_5_io_outHeadFlit_priorityLevel ),
       .io_result( CMeshDOR_5_io_result ),
       .io_vcsAvailable_4( CMeshDOR_5_io_vcsAvailable_4 ),
       .io_vcsAvailable_3( CMeshDOR_5_io_vcsAvailable_3 ),
       .io_vcsAvailable_2( CMeshDOR_5_io_vcsAvailable_2 ),
       .io_vcsAvailable_1( CMeshDOR_5_io_vcsAvailable_1 ),
       .io_vcsAvailable_0( CMeshDOR_5_io_vcsAvailable_0 )
  );
  VCRouterStateManagement VCRouterStateManagement_5(.clk(clk), .reset(reset),
       .io_inputBufferValid( RouterBuffer_5_io_deq_valid ),
       .io_routingComplete( R925 ),
       .io_inputBufferIsTail( T916 ),
       .io_vcAllocGranted( vcAllocator_io_resources_5_valid ),
       .io_swAllocGranted( T896 ),
       .io_creditsAvail( T877 ),
       .io_outputReady( T864 ),
       .io_currentState( VCRouterStateManagement_5_io_currentState )
  );
  ReplaceVCPort ReplaceVCPort_5(
       .io_oldFlit_x( T862 ),
       .io_newVCPort( T3140 ),
       .io_newFlit_x( ReplaceVCPort_5_io_newFlit_x )
  );
  Flit2FlitBundle Flit2FlitBundle_5(
       .io_inFlit_x( T856 )
       //.io_outHead_packetID(  )
       //.io_outHead_isTail(  )
       //.io_outHead_vcPort(  )
       //.io_outHead_packetType(  )
       //.io_outHead_destination_2(  )
       //.io_outHead_destination_1(  )
       //.io_outHead_destination_0(  )
       //.io_outHead_priorityLevel(  )
       //.io_outBody_packetID(  )
       //.io_outBody_isTail(  )
       //.io_outBody_vcPort(  )
       //.io_outBody_flitID(  )
       //.io_outBody_payload(  )
  );
  CreditGen CreditGen_6(
       .io_outCredit_grant( CreditGen_6_io_outCredit_grant ),
       .io_inGrant( T846 )
  );
  RouterRegFile RouterRegFile_6(.clk(clk), .reset(reset),
       .io_writeData( T844 ),
       .io_writeEnable( T841 ),
       //.io_full(  )
       .io_readData( RouterRegFile_6_io_readData ),
       .io_readValid( RouterRegFile_6_io_readValid ),
       .io_readIncrement( T828 ),
       .io_writePipelineReg_2( RouterRegFile_6_io_readPipelineReg_1 ),
       .io_writePipelineReg_1( RouterRegFile_6_io_readPipelineReg_0 ),
       .io_writePipelineReg_0( T3139 ),
       .io_wePipelineReg_2( T817 ),
       .io_wePipelineReg_1( T814 ),
       .io_wePipelineReg_0( T812 ),
       //.io_readPipelineReg_2(  )
       .io_readPipelineReg_1( RouterRegFile_6_io_readPipelineReg_1 ),
       .io_readPipelineReg_0( RouterRegFile_6_io_readPipelineReg_0 ),
       //.io_rvPipelineReg_2(  )
       .io_rvPipelineReg_1( RouterRegFile_6_io_rvPipelineReg_1 ),
       .io_rvPipelineReg_0( RouterRegFile_6_io_rvPipelineReg_0 )
  );
  RouterBuffer RouterBuffer_6(.clk(clk), .reset(reset),
       .io_enq_ready( RouterBuffer_6_io_enq_ready ),
       .io_enq_valid( T811 ),
       .io_enq_bits_x( io_inChannels_3_flit_x ),
       .io_deq_ready( T792 ),
       .io_deq_valid( RouterBuffer_6_io_deq_valid ),
       .io_deq_bits_x( RouterBuffer_6_io_deq_bits_x )
  );
  CMeshDOR_2 CMeshDOR_6(
       .io_inHeadFlit_packetID( T791 ),
       .io_inHeadFlit_isTail( T790 ),
       .io_inHeadFlit_vcPort( T789 ),
       .io_inHeadFlit_packetType( T788 ),
       .io_inHeadFlit_destination_2( T787 ),
       .io_inHeadFlit_destination_1( T786 ),
       .io_inHeadFlit_destination_0( T785 ),
       .io_inHeadFlit_priorityLevel( T782 ),
       .io_outHeadFlit_packetID( CMeshDOR_6_io_outHeadFlit_packetID ),
       .io_outHeadFlit_isTail( CMeshDOR_6_io_outHeadFlit_isTail ),
       .io_outHeadFlit_vcPort( CMeshDOR_6_io_outHeadFlit_vcPort ),
       .io_outHeadFlit_packetType( CMeshDOR_6_io_outHeadFlit_packetType ),
       .io_outHeadFlit_destination_2( CMeshDOR_6_io_outHeadFlit_destination_2 ),
       .io_outHeadFlit_destination_1( CMeshDOR_6_io_outHeadFlit_destination_1 ),
       .io_outHeadFlit_destination_0( CMeshDOR_6_io_outHeadFlit_destination_0 ),
       .io_outHeadFlit_priorityLevel( CMeshDOR_6_io_outHeadFlit_priorityLevel ),
       .io_result( CMeshDOR_6_io_result ),
       .io_vcsAvailable_4( CMeshDOR_6_io_vcsAvailable_4 ),
       .io_vcsAvailable_3( CMeshDOR_6_io_vcsAvailable_3 ),
       .io_vcsAvailable_2( CMeshDOR_6_io_vcsAvailable_2 ),
       .io_vcsAvailable_1( CMeshDOR_6_io_vcsAvailable_1 ),
       .io_vcsAvailable_0( CMeshDOR_6_io_vcsAvailable_0 )
  );
  VCRouterStateManagement VCRouterStateManagement_6(.clk(clk), .reset(reset),
       .io_inputBufferValid( RouterBuffer_6_io_deq_valid ),
       .io_routingComplete( R781 ),
       .io_inputBufferIsTail( T772 ),
       .io_vcAllocGranted( vcAllocator_io_resources_6_valid ),
       .io_swAllocGranted( T752 ),
       .io_creditsAvail( T733 ),
       .io_outputReady( T720 ),
       .io_currentState( VCRouterStateManagement_6_io_currentState )
  );
  ReplaceVCPort ReplaceVCPort_6(
       .io_oldFlit_x( T718 ),
       .io_newVCPort( T3133 ),
       .io_newFlit_x( ReplaceVCPort_6_io_newFlit_x )
  );
  Flit2FlitBundle Flit2FlitBundle_6(
       .io_inFlit_x( T712 )
       //.io_outHead_packetID(  )
       //.io_outHead_isTail(  )
       //.io_outHead_vcPort(  )
       //.io_outHead_packetType(  )
       //.io_outHead_destination_2(  )
       //.io_outHead_destination_1(  )
       //.io_outHead_destination_0(  )
       //.io_outHead_priorityLevel(  )
       //.io_outBody_packetID(  )
       //.io_outBody_isTail(  )
       //.io_outBody_vcPort(  )
       //.io_outBody_flitID(  )
       //.io_outBody_payload(  )
  );
  CreditGen CreditGen_7(
       .io_outCredit_grant( CreditGen_7_io_outCredit_grant ),
       .io_inGrant( T702 )
  );
  RouterRegFile RouterRegFile_7(.clk(clk), .reset(reset),
       .io_writeData( T700 ),
       .io_writeEnable( T697 ),
       //.io_full(  )
       .io_readData( RouterRegFile_7_io_readData ),
       .io_readValid( RouterRegFile_7_io_readValid ),
       .io_readIncrement( T684 ),
       .io_writePipelineReg_2( RouterRegFile_7_io_readPipelineReg_1 ),
       .io_writePipelineReg_1( RouterRegFile_7_io_readPipelineReg_0 ),
       .io_writePipelineReg_0( T3132 ),
       .io_wePipelineReg_2( T673 ),
       .io_wePipelineReg_1( T670 ),
       .io_wePipelineReg_0( T668 ),
       //.io_readPipelineReg_2(  )
       .io_readPipelineReg_1( RouterRegFile_7_io_readPipelineReg_1 ),
       .io_readPipelineReg_0( RouterRegFile_7_io_readPipelineReg_0 ),
       //.io_rvPipelineReg_2(  )
       .io_rvPipelineReg_1( RouterRegFile_7_io_rvPipelineReg_1 ),
       .io_rvPipelineReg_0( RouterRegFile_7_io_rvPipelineReg_0 )
  );
  RouterBuffer RouterBuffer_7(.clk(clk), .reset(reset),
       .io_enq_ready( RouterBuffer_7_io_enq_ready ),
       .io_enq_valid( T667 ),
       .io_enq_bits_x( io_inChannels_3_flit_x ),
       .io_deq_ready( T648 ),
       .io_deq_valid( RouterBuffer_7_io_deq_valid ),
       .io_deq_bits_x( RouterBuffer_7_io_deq_bits_x )
  );
  CMeshDOR_2 CMeshDOR_7(
       .io_inHeadFlit_packetID( T647 ),
       .io_inHeadFlit_isTail( T646 ),
       .io_inHeadFlit_vcPort( T645 ),
       .io_inHeadFlit_packetType( T644 ),
       .io_inHeadFlit_destination_2( T643 ),
       .io_inHeadFlit_destination_1( T642 ),
       .io_inHeadFlit_destination_0( T641 ),
       .io_inHeadFlit_priorityLevel( T638 ),
       .io_outHeadFlit_packetID( CMeshDOR_7_io_outHeadFlit_packetID ),
       .io_outHeadFlit_isTail( CMeshDOR_7_io_outHeadFlit_isTail ),
       .io_outHeadFlit_vcPort( CMeshDOR_7_io_outHeadFlit_vcPort ),
       .io_outHeadFlit_packetType( CMeshDOR_7_io_outHeadFlit_packetType ),
       .io_outHeadFlit_destination_2( CMeshDOR_7_io_outHeadFlit_destination_2 ),
       .io_outHeadFlit_destination_1( CMeshDOR_7_io_outHeadFlit_destination_1 ),
       .io_outHeadFlit_destination_0( CMeshDOR_7_io_outHeadFlit_destination_0 ),
       .io_outHeadFlit_priorityLevel( CMeshDOR_7_io_outHeadFlit_priorityLevel ),
       .io_result( CMeshDOR_7_io_result ),
       .io_vcsAvailable_4( CMeshDOR_7_io_vcsAvailable_4 ),
       .io_vcsAvailable_3( CMeshDOR_7_io_vcsAvailable_3 ),
       .io_vcsAvailable_2( CMeshDOR_7_io_vcsAvailable_2 ),
       .io_vcsAvailable_1( CMeshDOR_7_io_vcsAvailable_1 ),
       .io_vcsAvailable_0( CMeshDOR_7_io_vcsAvailable_0 )
  );
  VCRouterStateManagement VCRouterStateManagement_7(.clk(clk), .reset(reset),
       .io_inputBufferValid( RouterBuffer_7_io_deq_valid ),
       .io_routingComplete( R637 ),
       .io_inputBufferIsTail( T628 ),
       .io_vcAllocGranted( vcAllocator_io_resources_7_valid ),
       .io_swAllocGranted( T608 ),
       .io_creditsAvail( T589 ),
       .io_outputReady( T576 ),
       .io_currentState( VCRouterStateManagement_7_io_currentState )
  );
  ReplaceVCPort ReplaceVCPort_7(
       .io_oldFlit_x( T574 ),
       .io_newVCPort( T3126 ),
       .io_newFlit_x( ReplaceVCPort_7_io_newFlit_x )
  );
  Flit2FlitBundle Flit2FlitBundle_7(
       .io_inFlit_x( T568 )
       //.io_outHead_packetID(  )
       //.io_outHead_isTail(  )
       //.io_outHead_vcPort(  )
       //.io_outHead_packetType(  )
       //.io_outHead_destination_2(  )
       //.io_outHead_destination_1(  )
       //.io_outHead_destination_0(  )
       //.io_outHead_priorityLevel(  )
       //.io_outBody_packetID(  )
       //.io_outBody_isTail(  )
       //.io_outBody_vcPort(  )
       //.io_outBody_flitID(  )
       //.io_outBody_payload(  )
  );
  CreditGen CreditGen_8(
       .io_outCredit_grant( CreditGen_8_io_outCredit_grant ),
       .io_inGrant( T558 )
  );
  RouterRegFile RouterRegFile_8(.clk(clk), .reset(reset),
       .io_writeData( T556 ),
       .io_writeEnable( T553 ),
       //.io_full(  )
       .io_readData( RouterRegFile_8_io_readData ),
       .io_readValid( RouterRegFile_8_io_readValid ),
       .io_readIncrement( T540 ),
       .io_writePipelineReg_2( RouterRegFile_8_io_readPipelineReg_1 ),
       .io_writePipelineReg_1( RouterRegFile_8_io_readPipelineReg_0 ),
       .io_writePipelineReg_0( T3125 ),
       .io_wePipelineReg_2( T529 ),
       .io_wePipelineReg_1( T526 ),
       .io_wePipelineReg_0( T524 ),
       //.io_readPipelineReg_2(  )
       .io_readPipelineReg_1( RouterRegFile_8_io_readPipelineReg_1 ),
       .io_readPipelineReg_0( RouterRegFile_8_io_readPipelineReg_0 ),
       //.io_rvPipelineReg_2(  )
       .io_rvPipelineReg_1( RouterRegFile_8_io_rvPipelineReg_1 ),
       .io_rvPipelineReg_0( RouterRegFile_8_io_rvPipelineReg_0 )
  );
  RouterBuffer RouterBuffer_8(.clk(clk), .reset(reset),
       .io_enq_ready( RouterBuffer_8_io_enq_ready ),
       .io_enq_valid( T523 ),
       .io_enq_bits_x( io_inChannels_4_flit_x ),
       .io_deq_ready( T504 ),
       .io_deq_valid( RouterBuffer_8_io_deq_valid ),
       .io_deq_bits_x( RouterBuffer_8_io_deq_bits_x )
  );
  CMeshDOR_2 CMeshDOR_8(
       .io_inHeadFlit_packetID( T503 ),
       .io_inHeadFlit_isTail( T502 ),
       .io_inHeadFlit_vcPort( T501 ),
       .io_inHeadFlit_packetType( T500 ),
       .io_inHeadFlit_destination_2( T499 ),
       .io_inHeadFlit_destination_1( T498 ),
       .io_inHeadFlit_destination_0( T497 ),
       .io_inHeadFlit_priorityLevel( T494 ),
       .io_outHeadFlit_packetID( CMeshDOR_8_io_outHeadFlit_packetID ),
       .io_outHeadFlit_isTail( CMeshDOR_8_io_outHeadFlit_isTail ),
       .io_outHeadFlit_vcPort( CMeshDOR_8_io_outHeadFlit_vcPort ),
       .io_outHeadFlit_packetType( CMeshDOR_8_io_outHeadFlit_packetType ),
       .io_outHeadFlit_destination_2( CMeshDOR_8_io_outHeadFlit_destination_2 ),
       .io_outHeadFlit_destination_1( CMeshDOR_8_io_outHeadFlit_destination_1 ),
       .io_outHeadFlit_destination_0( CMeshDOR_8_io_outHeadFlit_destination_0 ),
       .io_outHeadFlit_priorityLevel( CMeshDOR_8_io_outHeadFlit_priorityLevel ),
       .io_result( CMeshDOR_8_io_result ),
       .io_vcsAvailable_4( CMeshDOR_8_io_vcsAvailable_4 ),
       .io_vcsAvailable_3( CMeshDOR_8_io_vcsAvailable_3 ),
       .io_vcsAvailable_2( CMeshDOR_8_io_vcsAvailable_2 ),
       .io_vcsAvailable_1( CMeshDOR_8_io_vcsAvailable_1 ),
       .io_vcsAvailable_0( CMeshDOR_8_io_vcsAvailable_0 )
  );
  VCRouterStateManagement VCRouterStateManagement_8(.clk(clk), .reset(reset),
       .io_inputBufferValid( RouterBuffer_8_io_deq_valid ),
       .io_routingComplete( R493 ),
       .io_inputBufferIsTail( T484 ),
       .io_vcAllocGranted( vcAllocator_io_resources_8_valid ),
       .io_swAllocGranted( T464 ),
       .io_creditsAvail( T445 ),
       .io_outputReady( T432 ),
       .io_currentState( VCRouterStateManagement_8_io_currentState )
  );
  ReplaceVCPort ReplaceVCPort_8(
       .io_oldFlit_x( T430 ),
       .io_newVCPort( T3119 ),
       .io_newFlit_x( ReplaceVCPort_8_io_newFlit_x )
  );
  Flit2FlitBundle Flit2FlitBundle_8(
       .io_inFlit_x( T424 )
       //.io_outHead_packetID(  )
       //.io_outHead_isTail(  )
       //.io_outHead_vcPort(  )
       //.io_outHead_packetType(  )
       //.io_outHead_destination_2(  )
       //.io_outHead_destination_1(  )
       //.io_outHead_destination_0(  )
       //.io_outHead_priorityLevel(  )
       //.io_outBody_packetID(  )
       //.io_outBody_isTail(  )
       //.io_outBody_vcPort(  )
       //.io_outBody_flitID(  )
       //.io_outBody_payload(  )
  );
  CreditGen CreditGen_9(
       .io_outCredit_grant( CreditGen_9_io_outCredit_grant ),
       .io_inGrant( T414 )
  );
  RouterRegFile RouterRegFile_9(.clk(clk), .reset(reset),
       .io_writeData( T412 ),
       .io_writeEnable( T409 ),
       //.io_full(  )
       .io_readData( RouterRegFile_9_io_readData ),
       .io_readValid( RouterRegFile_9_io_readValid ),
       .io_readIncrement( T396 ),
       .io_writePipelineReg_2( RouterRegFile_9_io_readPipelineReg_1 ),
       .io_writePipelineReg_1( RouterRegFile_9_io_readPipelineReg_0 ),
       .io_writePipelineReg_0( T3118 ),
       .io_wePipelineReg_2( T385 ),
       .io_wePipelineReg_1( T382 ),
       .io_wePipelineReg_0( T380 ),
       //.io_readPipelineReg_2(  )
       .io_readPipelineReg_1( RouterRegFile_9_io_readPipelineReg_1 ),
       .io_readPipelineReg_0( RouterRegFile_9_io_readPipelineReg_0 ),
       //.io_rvPipelineReg_2(  )
       .io_rvPipelineReg_1( RouterRegFile_9_io_rvPipelineReg_1 ),
       .io_rvPipelineReg_0( RouterRegFile_9_io_rvPipelineReg_0 )
  );
  RouterBuffer RouterBuffer_9(.clk(clk), .reset(reset),
       .io_enq_ready( RouterBuffer_9_io_enq_ready ),
       .io_enq_valid( T379 ),
       .io_enq_bits_x( io_inChannels_4_flit_x ),
       .io_deq_ready( T360 ),
       .io_deq_valid( RouterBuffer_9_io_deq_valid ),
       .io_deq_bits_x( RouterBuffer_9_io_deq_bits_x )
  );
  CMeshDOR_2 CMeshDOR_9(
       .io_inHeadFlit_packetID( T359 ),
       .io_inHeadFlit_isTail( T358 ),
       .io_inHeadFlit_vcPort( T357 ),
       .io_inHeadFlit_packetType( T356 ),
       .io_inHeadFlit_destination_2( T355 ),
       .io_inHeadFlit_destination_1( T354 ),
       .io_inHeadFlit_destination_0( T353 ),
       .io_inHeadFlit_priorityLevel( T350 ),
       .io_outHeadFlit_packetID( CMeshDOR_9_io_outHeadFlit_packetID ),
       .io_outHeadFlit_isTail( CMeshDOR_9_io_outHeadFlit_isTail ),
       .io_outHeadFlit_vcPort( CMeshDOR_9_io_outHeadFlit_vcPort ),
       .io_outHeadFlit_packetType( CMeshDOR_9_io_outHeadFlit_packetType ),
       .io_outHeadFlit_destination_2( CMeshDOR_9_io_outHeadFlit_destination_2 ),
       .io_outHeadFlit_destination_1( CMeshDOR_9_io_outHeadFlit_destination_1 ),
       .io_outHeadFlit_destination_0( CMeshDOR_9_io_outHeadFlit_destination_0 ),
       .io_outHeadFlit_priorityLevel( CMeshDOR_9_io_outHeadFlit_priorityLevel ),
       .io_result( CMeshDOR_9_io_result ),
       .io_vcsAvailable_4( CMeshDOR_9_io_vcsAvailable_4 ),
       .io_vcsAvailable_3( CMeshDOR_9_io_vcsAvailable_3 ),
       .io_vcsAvailable_2( CMeshDOR_9_io_vcsAvailable_2 ),
       .io_vcsAvailable_1( CMeshDOR_9_io_vcsAvailable_1 ),
       .io_vcsAvailable_0( CMeshDOR_9_io_vcsAvailable_0 )
  );
  VCRouterStateManagement VCRouterStateManagement_9(.clk(clk), .reset(reset),
       .io_inputBufferValid( RouterBuffer_9_io_deq_valid ),
       .io_routingComplete( R349 ),
       .io_inputBufferIsTail( T340 ),
       .io_vcAllocGranted( vcAllocator_io_resources_9_valid ),
       .io_swAllocGranted( T320 ),
       .io_creditsAvail( T301 ),
       .io_outputReady( T288 ),
       .io_currentState( VCRouterStateManagement_9_io_currentState )
  );
  ReplaceVCPort ReplaceVCPort_9(
       .io_oldFlit_x( T286 ),
       .io_newVCPort( T3112 ),
       .io_newFlit_x( ReplaceVCPort_9_io_newFlit_x )
  );
  Flit2FlitBundle Flit2FlitBundle_9(
       .io_inFlit_x( T280 )
       //.io_outHead_packetID(  )
       //.io_outHead_isTail(  )
       //.io_outHead_vcPort(  )
       //.io_outHead_packetType(  )
       //.io_outHead_destination_2(  )
       //.io_outHead_destination_1(  )
       //.io_outHead_destination_0(  )
       //.io_outHead_priorityLevel(  )
       //.io_outBody_packetID(  )
       //.io_outBody_isTail(  )
       //.io_outBody_vcPort(  )
       //.io_outBody_flitID(  )
       //.io_outBody_payload(  )
  );
  CreditCon CreditCon(.clk(clk), .reset(reset),
       .io_inCredit_grant( io_outChannels_0_credit_0_grant ),
       .io_inConsume( T278 ),
       .io_outCredit( CreditCon_io_outCredit )
       //.io_almostOut(  )
  );
  CreditCon CreditCon_1(.clk(clk), .reset(reset),
       .io_inCredit_grant( io_outChannels_0_credit_1_grant ),
       .io_inConsume( T268 ),
       .io_outCredit( CreditCon_1_io_outCredit )
       //.io_almostOut(  )
  );
  MuxN_1 MuxN(
       //.io_ins_1(  )
       //.io_ins_0(  )
       //.io_sel(  )
       //.io_out(  )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign MuxN.io_ins_1 = {1{1'b0}};
    assign MuxN.io_ins_0 = {1{1'b0}};
    assign MuxN.io_sel = {1{1'b0}};
// synthesis translate_on
`endif
  CreditCon CreditCon_2(.clk(clk), .reset(reset),
       .io_inCredit_grant( io_outChannels_1_credit_0_grant ),
       .io_inConsume( T266 ),
       .io_outCredit( CreditCon_2_io_outCredit )
       //.io_almostOut(  )
  );
  CreditCon CreditCon_3(.clk(clk), .reset(reset),
       .io_inCredit_grant( io_outChannels_1_credit_1_grant ),
       .io_inConsume( T256 ),
       .io_outCredit( CreditCon_3_io_outCredit )
       //.io_almostOut(  )
  );
  MuxN_1 MuxN_1(
       //.io_ins_1(  )
       //.io_ins_0(  )
       //.io_sel(  )
       //.io_out(  )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign MuxN_1.io_ins_1 = {1{1'b0}};
    assign MuxN_1.io_ins_0 = {1{1'b0}};
    assign MuxN_1.io_sel = {1{1'b0}};
// synthesis translate_on
`endif
  CreditCon CreditCon_4(.clk(clk), .reset(reset),
       .io_inCredit_grant( io_outChannels_2_credit_0_grant ),
       .io_inConsume( T254 ),
       .io_outCredit( CreditCon_4_io_outCredit )
       //.io_almostOut(  )
  );
  CreditCon CreditCon_5(.clk(clk), .reset(reset),
       .io_inCredit_grant( io_outChannels_2_credit_1_grant ),
       .io_inConsume( T244 ),
       .io_outCredit( CreditCon_5_io_outCredit )
       //.io_almostOut(  )
  );
  MuxN_1 MuxN_2(
       //.io_ins_1(  )
       //.io_ins_0(  )
       //.io_sel(  )
       //.io_out(  )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign MuxN_2.io_ins_1 = {1{1'b0}};
    assign MuxN_2.io_ins_0 = {1{1'b0}};
    assign MuxN_2.io_sel = {1{1'b0}};
// synthesis translate_on
`endif
  CreditCon CreditCon_6(.clk(clk), .reset(reset),
       .io_inCredit_grant( io_outChannels_3_credit_0_grant ),
       .io_inConsume( T242 ),
       .io_outCredit( CreditCon_6_io_outCredit )
       //.io_almostOut(  )
  );
  CreditCon CreditCon_7(.clk(clk), .reset(reset),
       .io_inCredit_grant( io_outChannels_3_credit_1_grant ),
       .io_inConsume( T232 ),
       .io_outCredit( CreditCon_7_io_outCredit )
       //.io_almostOut(  )
  );
  MuxN_1 MuxN_3(
       //.io_ins_1(  )
       //.io_ins_0(  )
       //.io_sel(  )
       //.io_out(  )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign MuxN_3.io_ins_1 = {1{1'b0}};
    assign MuxN_3.io_ins_0 = {1{1'b0}};
    assign MuxN_3.io_sel = {1{1'b0}};
// synthesis translate_on
`endif
  CreditCon CreditCon_8(.clk(clk), .reset(reset),
       .io_inCredit_grant( io_outChannels_4_credit_0_grant ),
       .io_inConsume( T230 ),
       .io_outCredit( CreditCon_8_io_outCredit )
       //.io_almostOut(  )
  );
  CreditCon CreditCon_9(.clk(clk), .reset(reset),
       .io_inCredit_grant( io_outChannels_4_credit_1_grant ),
       .io_inConsume( T220 ),
       .io_outCredit( CreditCon_9_io_outCredit )
       //.io_almostOut(  )
  );
  MuxN_1 MuxN_4(
       //.io_ins_1(  )
       //.io_ins_0(  )
       //.io_sel(  )
       //.io_out(  )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign MuxN_4.io_ins_1 = {1{1'b0}};
    assign MuxN_4.io_ins_0 = {1{1'b0}};
    assign MuxN_4.io_sel = {1{1'b0}};
// synthesis translate_on
`endif

  always @(posedge clk) begin
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T215 <= 1'b1;
  if(!T216 && T215 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "SimpleVCRouter: Flit with VC port/*? in < (class OpenSoC.SimpleVCRouter)>*/ Chisel.UInt(width=1, connect to 1 inputs: ([Chisel.Mux] in OpenSoC.SimpleVCRouter)) attempting to write to VC 0");
    $finish;
  end
// synthesis translate_on
`endif
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T198 <= 1'b1;
  if(!T199 && T198 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "SimpleVCRouter:Vector(2, 0) Insufficent space in input buffer - Credit Ready asserted when Routing In Buffer not ready inputPort= 0 curVC = 0");
    $finish;
  end
// synthesis translate_on
`endif
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T193 <= 1'b1;
  if(!T194 && T193 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "SimpleVCRouter: Flit with VC port/*? in < (class OpenSoC.SimpleVCRouter)>*/ Chisel.UInt(width=1, connect to 1 inputs: ([Chisel.Mux] in OpenSoC.SimpleVCRouter)) attempting to write to VC 1");
    $finish;
  end
// synthesis translate_on
`endif
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T176 <= 1'b1;
  if(!T177 && T176 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "SimpleVCRouter:Vector(2, 0) Insufficent space in input buffer - Credit Ready asserted when Routing In Buffer not ready inputPort= 0 curVC = 1");
    $finish;
  end
// synthesis translate_on
`endif
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T171 <= 1'b1;
  if(!T172 && T171 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "SimpleVCRouter: Flit with VC port/*? in < (class OpenSoC.SimpleVCRouter)>*/ Chisel.UInt(width=1, connect to 1 inputs: ([Chisel.Mux] in OpenSoC.SimpleVCRouter)) attempting to write to VC 0");
    $finish;
  end
// synthesis translate_on
`endif
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T154 <= 1'b1;
  if(!T155 && T154 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "SimpleVCRouter:Vector(2, 0) Insufficent space in input buffer - Credit Ready asserted when Routing In Buffer not ready inputPort= 1 curVC = 0");
    $finish;
  end
// synthesis translate_on
`endif
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T149 <= 1'b1;
  if(!T150 && T149 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "SimpleVCRouter: Flit with VC port/*? in < (class OpenSoC.SimpleVCRouter)>*/ Chisel.UInt(width=1, connect to 1 inputs: ([Chisel.Mux] in OpenSoC.SimpleVCRouter)) attempting to write to VC 1");
    $finish;
  end
// synthesis translate_on
`endif
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T132 <= 1'b1;
  if(!T133 && T132 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "SimpleVCRouter:Vector(2, 0) Insufficent space in input buffer - Credit Ready asserted when Routing In Buffer not ready inputPort= 1 curVC = 1");
    $finish;
  end
// synthesis translate_on
`endif
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T127 <= 1'b1;
  if(!T128 && T127 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "SimpleVCRouter: Flit with VC port/*? in < (class OpenSoC.SimpleVCRouter)>*/ Chisel.UInt(width=1, connect to 1 inputs: ([Chisel.Mux] in OpenSoC.SimpleVCRouter)) attempting to write to VC 0");
    $finish;
  end
// synthesis translate_on
`endif
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T110 <= 1'b1;
  if(!T111 && T110 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "SimpleVCRouter:Vector(2, 0) Insufficent space in input buffer - Credit Ready asserted when Routing In Buffer not ready inputPort= 2 curVC = 0");
    $finish;
  end
// synthesis translate_on
`endif
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T105 <= 1'b1;
  if(!T106 && T105 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "SimpleVCRouter: Flit with VC port/*? in < (class OpenSoC.SimpleVCRouter)>*/ Chisel.UInt(width=1, connect to 1 inputs: ([Chisel.Mux] in OpenSoC.SimpleVCRouter)) attempting to write to VC 1");
    $finish;
  end
// synthesis translate_on
`endif
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T88 <= 1'b1;
  if(!T89 && T88 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "SimpleVCRouter:Vector(2, 0) Insufficent space in input buffer - Credit Ready asserted when Routing In Buffer not ready inputPort= 2 curVC = 1");
    $finish;
  end
// synthesis translate_on
`endif
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T83 <= 1'b1;
  if(!T84 && T83 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "SimpleVCRouter: Flit with VC port/*? in < (class OpenSoC.SimpleVCRouter)>*/ Chisel.UInt(width=1, connect to 1 inputs: ([Chisel.Mux] in OpenSoC.SimpleVCRouter)) attempting to write to VC 0");
    $finish;
  end
// synthesis translate_on
`endif
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T66 <= 1'b1;
  if(!T67 && T66 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "SimpleVCRouter:Vector(2, 0) Insufficent space in input buffer - Credit Ready asserted when Routing In Buffer not ready inputPort= 3 curVC = 0");
    $finish;
  end
// synthesis translate_on
`endif
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T61 <= 1'b1;
  if(!T62 && T61 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "SimpleVCRouter: Flit with VC port/*? in < (class OpenSoC.SimpleVCRouter)>*/ Chisel.UInt(width=1, connect to 1 inputs: ([Chisel.Mux] in OpenSoC.SimpleVCRouter)) attempting to write to VC 1");
    $finish;
  end
// synthesis translate_on
`endif
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T44 <= 1'b1;
  if(!T45 && T44 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "SimpleVCRouter:Vector(2, 0) Insufficent space in input buffer - Credit Ready asserted when Routing In Buffer not ready inputPort= 3 curVC = 1");
    $finish;
  end
// synthesis translate_on
`endif
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T39 <= 1'b1;
  if(!T40 && T39 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "SimpleVCRouter: Flit with VC port/*? in < (class OpenSoC.SimpleVCRouter)>*/ Chisel.UInt(width=1, connect to 1 inputs: ([Chisel.Mux] in OpenSoC.SimpleVCRouter)) attempting to write to VC 0");
    $finish;
  end
// synthesis translate_on
`endif
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T22 <= 1'b1;
  if(!T23 && T22 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "SimpleVCRouter:Vector(2, 0) Insufficent space in input buffer - Credit Ready asserted when Routing In Buffer not ready inputPort= 4 curVC = 0");
    $finish;
  end
// synthesis translate_on
`endif
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T17 <= 1'b1;
  if(!T18 && T17 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "SimpleVCRouter: Flit with VC port/*? in < (class OpenSoC.SimpleVCRouter)>*/ Chisel.UInt(width=1, connect to 1 inputs: ([Chisel.Mux] in OpenSoC.SimpleVCRouter)) attempting to write to VC 1");
    $finish;
  end
// synthesis translate_on
`endif
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T0 <= 1'b1;
  if(!T1 && T0 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "SimpleVCRouter:Vector(2, 0) Insufficent space in input buffer - Credit Ready asserted when Routing In Buffer not ready inputPort= 4 curVC = 1");
    $finish;
  end
// synthesis translate_on
`endif
    if(reset) begin
      R282 <= 55'h0;
    end else if(T284) begin
      R282 <= T3114;
    end
    if(reset) begin
      R295 <= 3'h0;
    end else begin
      R295 <= CMeshDOR_9_io_result;
    end
    if(reset) begin
      R349 <= 1'h0;
    end else begin
      R349 <= RouterBuffer_9_io_deq_valid;
    end
    if(reset) begin
      R426 <= 55'h0;
    end else if(T428) begin
      R426 <= T3121;
    end
    if(reset) begin
      R439 <= 3'h0;
    end else begin
      R439 <= CMeshDOR_8_io_result;
    end
    if(reset) begin
      R493 <= 1'h0;
    end else begin
      R493 <= RouterBuffer_8_io_deq_valid;
    end
    if(reset) begin
      R570 <= 55'h0;
    end else if(T572) begin
      R570 <= T3128;
    end
    if(reset) begin
      R583 <= 3'h0;
    end else begin
      R583 <= CMeshDOR_7_io_result;
    end
    if(reset) begin
      R637 <= 1'h0;
    end else begin
      R637 <= RouterBuffer_7_io_deq_valid;
    end
    if(reset) begin
      R714 <= 55'h0;
    end else if(T716) begin
      R714 <= T3135;
    end
    if(reset) begin
      R727 <= 3'h0;
    end else begin
      R727 <= CMeshDOR_6_io_result;
    end
    if(reset) begin
      R781 <= 1'h0;
    end else begin
      R781 <= RouterBuffer_6_io_deq_valid;
    end
    if(reset) begin
      R858 <= 55'h0;
    end else if(T860) begin
      R858 <= T3142;
    end
    if(reset) begin
      R871 <= 3'h0;
    end else begin
      R871 <= CMeshDOR_5_io_result;
    end
    if(reset) begin
      R925 <= 1'h0;
    end else begin
      R925 <= RouterBuffer_5_io_deq_valid;
    end
    if(reset) begin
      R1002 <= 55'h0;
    end else if(T1004) begin
      R1002 <= T3149;
    end
    if(reset) begin
      R1015 <= 3'h0;
    end else begin
      R1015 <= CMeshDOR_4_io_result;
    end
    if(reset) begin
      R1069 <= 1'h0;
    end else begin
      R1069 <= RouterBuffer_4_io_deq_valid;
    end
    if(reset) begin
      R1146 <= 55'h0;
    end else if(T1148) begin
      R1146 <= T3156;
    end
    if(reset) begin
      R1159 <= 3'h0;
    end else begin
      R1159 <= CMeshDOR_3_io_result;
    end
    if(reset) begin
      R1213 <= 1'h0;
    end else begin
      R1213 <= RouterBuffer_3_io_deq_valid;
    end
    if(reset) begin
      R1290 <= 55'h0;
    end else if(T1292) begin
      R1290 <= T3163;
    end
    if(reset) begin
      R1303 <= 3'h0;
    end else begin
      R1303 <= CMeshDOR_2_io_result;
    end
    if(reset) begin
      R1357 <= 1'h0;
    end else begin
      R1357 <= RouterBuffer_2_io_deq_valid;
    end
    if(reset) begin
      R1434 <= 55'h0;
    end else if(T1436) begin
      R1434 <= T3170;
    end
    if(reset) begin
      R1447 <= 3'h0;
    end else begin
      R1447 <= CMeshDOR_1_io_result;
    end
    if(reset) begin
      R1501 <= 1'h0;
    end else begin
      R1501 <= RouterBuffer_1_io_deq_valid;
    end
    if(reset) begin
      R1578 <= 55'h0;
    end else if(T1580) begin
      R1578 <= T3177;
    end
    if(reset) begin
      R1591 <= 3'h0;
    end else begin
      R1591 <= CMeshDOR_io_result;
    end
    if(reset) begin
      R1645 <= 1'h0;
    end else begin
      R1645 <= RouterBuffer_io_deq_valid;
    end
    validVCs_0_0 <= CMeshDOR_io_vcsAvailable_0;
    R2176 <= T2177;
    R2181 <= T2182;
    validVCs_0_1 <= CMeshDOR_io_vcsAvailable_1;
    R2186 <= T2187;
    R2191 <= T2192;
    validVCs_0_2 <= CMeshDOR_io_vcsAvailable_2;
    R2196 <= T2197;
    R2201 <= T2202;
    validVCs_0_3 <= CMeshDOR_io_vcsAvailable_3;
    R2206 <= T2207;
    R2211 <= T2212;
    validVCs_0_4 <= CMeshDOR_io_vcsAvailable_4;
    R2216 <= T2217;
    R2221 <= T2222;
    validVCs_1_0 <= CMeshDOR_1_io_vcsAvailable_0;
    R2226 <= T2227;
    R2231 <= T2232;
    validVCs_1_1 <= CMeshDOR_1_io_vcsAvailable_1;
    R2236 <= T2237;
    R2241 <= T2242;
    validVCs_1_2 <= CMeshDOR_1_io_vcsAvailable_2;
    R2246 <= T2247;
    R2251 <= T2252;
    validVCs_1_3 <= CMeshDOR_1_io_vcsAvailable_3;
    R2256 <= T2257;
    R2261 <= T2262;
    validVCs_1_4 <= CMeshDOR_1_io_vcsAvailable_4;
    R2266 <= T2267;
    R2271 <= T2272;
    validVCs_2_0 <= CMeshDOR_2_io_vcsAvailable_0;
    R2276 <= T2277;
    R2281 <= T2282;
    validVCs_2_1 <= CMeshDOR_2_io_vcsAvailable_1;
    R2286 <= T2287;
    R2291 <= T2292;
    validVCs_2_2 <= CMeshDOR_2_io_vcsAvailable_2;
    R2296 <= T2297;
    R2301 <= T2302;
    validVCs_2_3 <= CMeshDOR_2_io_vcsAvailable_3;
    R2306 <= T2307;
    R2311 <= T2312;
    validVCs_2_4 <= CMeshDOR_2_io_vcsAvailable_4;
    R2316 <= T2317;
    R2321 <= T2322;
    validVCs_3_0 <= CMeshDOR_3_io_vcsAvailable_0;
    R2326 <= T2327;
    R2331 <= T2332;
    validVCs_3_1 <= CMeshDOR_3_io_vcsAvailable_1;
    R2336 <= T2337;
    R2341 <= T2342;
    validVCs_3_2 <= CMeshDOR_3_io_vcsAvailable_2;
    R2346 <= T2347;
    R2351 <= T2352;
    validVCs_3_3 <= CMeshDOR_3_io_vcsAvailable_3;
    R2356 <= T2357;
    R2361 <= T2362;
    validVCs_3_4 <= CMeshDOR_3_io_vcsAvailable_4;
    R2366 <= T2367;
    R2371 <= T2372;
    validVCs_4_0 <= CMeshDOR_4_io_vcsAvailable_0;
    R2376 <= T2377;
    R2381 <= T2382;
    validVCs_4_1 <= CMeshDOR_4_io_vcsAvailable_1;
    R2386 <= T2387;
    R2391 <= T2392;
    validVCs_4_2 <= CMeshDOR_4_io_vcsAvailable_2;
    R2396 <= T2397;
    R2401 <= T2402;
    validVCs_4_3 <= CMeshDOR_4_io_vcsAvailable_3;
    R2406 <= T2407;
    R2411 <= T2412;
    validVCs_4_4 <= CMeshDOR_4_io_vcsAvailable_4;
    R2416 <= T2417;
    R2421 <= T2422;
    validVCs_5_0 <= CMeshDOR_5_io_vcsAvailable_0;
    R2426 <= T2427;
    R2431 <= T2432;
    validVCs_5_1 <= CMeshDOR_5_io_vcsAvailable_1;
    R2436 <= T2437;
    R2441 <= T2442;
    validVCs_5_2 <= CMeshDOR_5_io_vcsAvailable_2;
    R2446 <= T2447;
    R2451 <= T2452;
    validVCs_5_3 <= CMeshDOR_5_io_vcsAvailable_3;
    R2456 <= T2457;
    R2461 <= T2462;
    validVCs_5_4 <= CMeshDOR_5_io_vcsAvailable_4;
    R2466 <= T2467;
    R2471 <= T2472;
    validVCs_6_0 <= CMeshDOR_6_io_vcsAvailable_0;
    R2476 <= T2477;
    R2481 <= T2482;
    validVCs_6_1 <= CMeshDOR_6_io_vcsAvailable_1;
    R2486 <= T2487;
    R2491 <= T2492;
    validVCs_6_2 <= CMeshDOR_6_io_vcsAvailable_2;
    R2496 <= T2497;
    R2501 <= T2502;
    validVCs_6_3 <= CMeshDOR_6_io_vcsAvailable_3;
    R2506 <= T2507;
    R2511 <= T2512;
    validVCs_6_4 <= CMeshDOR_6_io_vcsAvailable_4;
    R2516 <= T2517;
    R2521 <= T2522;
    validVCs_7_0 <= CMeshDOR_7_io_vcsAvailable_0;
    R2526 <= T2527;
    R2531 <= T2532;
    validVCs_7_1 <= CMeshDOR_7_io_vcsAvailable_1;
    R2536 <= T2537;
    R2541 <= T2542;
    validVCs_7_2 <= CMeshDOR_7_io_vcsAvailable_2;
    R2546 <= T2547;
    R2551 <= T2552;
    validVCs_7_3 <= CMeshDOR_7_io_vcsAvailable_3;
    R2556 <= T2557;
    R2561 <= T2562;
    validVCs_7_4 <= CMeshDOR_7_io_vcsAvailable_4;
    R2566 <= T2567;
    R2571 <= T2572;
    validVCs_8_0 <= CMeshDOR_8_io_vcsAvailable_0;
    R2576 <= T2577;
    R2581 <= T2582;
    validVCs_8_1 <= CMeshDOR_8_io_vcsAvailable_1;
    R2586 <= T2587;
    R2591 <= T2592;
    validVCs_8_2 <= CMeshDOR_8_io_vcsAvailable_2;
    R2596 <= T2597;
    R2601 <= T2602;
    validVCs_8_3 <= CMeshDOR_8_io_vcsAvailable_3;
    R2606 <= T2607;
    R2611 <= T2612;
    validVCs_8_4 <= CMeshDOR_8_io_vcsAvailable_4;
    R2616 <= T2617;
    R2621 <= T2622;
    validVCs_9_0 <= CMeshDOR_9_io_vcsAvailable_0;
    R2626 <= T2627;
    R2631 <= T2632;
    validVCs_9_1 <= CMeshDOR_9_io_vcsAvailable_1;
    R2636 <= T2637;
    R2641 <= T2642;
    validVCs_9_2 <= CMeshDOR_9_io_vcsAvailable_2;
    R2646 <= T2647;
    R2651 <= T2652;
    validVCs_9_3 <= CMeshDOR_9_io_vcsAvailable_3;
    R2656 <= T2657;
    R2661 <= T2662;
    validVCs_9_4 <= CMeshDOR_9_io_vcsAvailable_4;
    R2666 <= T2667;
    R2671 <= T2672;
    if(reset) begin
      R2675 <= 3'h0;
    end else if(T1670) begin
      R2675 <= T2677;
    end
    if(reset) begin
      R2683 <= 8'h0;
    end else begin
      R2683 <= T2684;
    end
    if(reset) begin
      R2688 <= 1'h1;
    end else begin
      R2688 <= T1692;
    end
    if(reset) begin
      R2689 <= 3'h0;
    end else if(T1526) begin
      R2689 <= T2691;
    end
    if(reset) begin
      R2697 <= 8'h0;
    end else begin
      R2697 <= T2698;
    end
    if(reset) begin
      R2702 <= 1'h1;
    end else begin
      R2702 <= T1548;
    end
    if(reset) begin
      R2703 <= 3'h0;
    end else if(T1382) begin
      R2703 <= T2705;
    end
    if(reset) begin
      R2711 <= 8'h0;
    end else begin
      R2711 <= T2712;
    end
    if(reset) begin
      R2716 <= 1'h1;
    end else begin
      R2716 <= T1404;
    end
    if(reset) begin
      R2717 <= 3'h0;
    end else if(T1238) begin
      R2717 <= T2719;
    end
    if(reset) begin
      R2725 <= 8'h0;
    end else begin
      R2725 <= T2726;
    end
    if(reset) begin
      R2730 <= 1'h1;
    end else begin
      R2730 <= T1260;
    end
    if(reset) begin
      R2731 <= 3'h0;
    end else if(T1094) begin
      R2731 <= T2733;
    end
    if(reset) begin
      R2739 <= 8'h0;
    end else begin
      R2739 <= T2740;
    end
    if(reset) begin
      R2744 <= 1'h1;
    end else begin
      R2744 <= T1116;
    end
    if(reset) begin
      R2745 <= 3'h0;
    end else if(T950) begin
      R2745 <= T2747;
    end
    if(reset) begin
      R2753 <= 8'h0;
    end else begin
      R2753 <= T2754;
    end
    if(reset) begin
      R2758 <= 1'h1;
    end else begin
      R2758 <= T972;
    end
    if(reset) begin
      R2759 <= 3'h0;
    end else if(T806) begin
      R2759 <= T2761;
    end
    if(reset) begin
      R2767 <= 8'h0;
    end else begin
      R2767 <= T2768;
    end
    if(reset) begin
      R2772 <= 1'h1;
    end else begin
      R2772 <= T828;
    end
    if(reset) begin
      R2773 <= 3'h0;
    end else if(T662) begin
      R2773 <= T2775;
    end
    if(reset) begin
      R2781 <= 8'h0;
    end else begin
      R2781 <= T2782;
    end
    if(reset) begin
      R2786 <= 1'h1;
    end else begin
      R2786 <= T684;
    end
    if(reset) begin
      R2787 <= 3'h0;
    end else if(T518) begin
      R2787 <= T2789;
    end
    if(reset) begin
      R2795 <= 8'h0;
    end else begin
      R2795 <= T2796;
    end
    if(reset) begin
      R2800 <= 1'h1;
    end else begin
      R2800 <= T540;
    end
    if(reset) begin
      R2801 <= 3'h0;
    end else if(T374) begin
      R2801 <= T2803;
    end
    if(reset) begin
      R2809 <= 8'h0;
    end else begin
      R2809 <= T2810;
    end
    if(reset) begin
      R2814 <= 1'h1;
    end else begin
      R2814 <= T396;
    end
    R3097 <= T2094;
    if(reset) begin
      R3098 <= T3099;
    end else begin
      R3098 <= switch_io_outPorts_0_x;
    end
    R3100 <= T2031;
    if(reset) begin
      R3101 <= T3102;
    end else begin
      R3101 <= switch_io_outPorts_1_x;
    end
    R3103 <= T1968;
    if(reset) begin
      R3104 <= T3105;
    end else begin
      R3104 <= switch_io_outPorts_2_x;
    end
    R3106 <= T1905;
    if(reset) begin
      R3107 <= T3108;
    end else begin
      R3107 <= switch_io_outPorts_3_x;
    end
    R3109 <= T1722;
    if(reset) begin
      R3110 <= T3111;
    end else begin
      R3110 <= switch_io_outPorts_4_x;
    end
  end
endmodule

module VCRouterWrapper_2(input clk, input reset,
    input [54:0] io_inChannels_4_flit_x,
    input  io_inChannels_4_flitValid,
    output io_inChannels_4_credit_1_grant,
    output io_inChannels_4_credit_0_grant,
    input [54:0] io_inChannels_3_flit_x,
    input  io_inChannels_3_flitValid,
    output io_inChannels_3_credit_1_grant,
    output io_inChannels_3_credit_0_grant,
    input [54:0] io_inChannels_2_flit_x,
    input  io_inChannels_2_flitValid,
    output io_inChannels_2_credit_1_grant,
    output io_inChannels_2_credit_0_grant,
    input [54:0] io_inChannels_1_flit_x,
    input  io_inChannels_1_flitValid,
    output io_inChannels_1_credit_1_grant,
    output io_inChannels_1_credit_0_grant,
    input [54:0] io_inChannels_0_flit_x,
    input  io_inChannels_0_flitValid,
    output io_inChannels_0_credit_1_grant,
    output io_inChannels_0_credit_0_grant,
    output[54:0] io_outChannels_4_flit_x,
    output io_outChannels_4_flitValid,
    input  io_outChannels_4_credit_1_grant,
    input  io_outChannels_4_credit_0_grant,
    output[54:0] io_outChannels_3_flit_x,
    output io_outChannels_3_flitValid,
    input  io_outChannels_3_credit_1_grant,
    input  io_outChannels_3_credit_0_grant,
    output[54:0] io_outChannels_2_flit_x,
    output io_outChannels_2_flitValid,
    input  io_outChannels_2_credit_1_grant,
    input  io_outChannels_2_credit_0_grant,
    output[54:0] io_outChannels_1_flit_x,
    output io_outChannels_1_flitValid,
    input  io_outChannels_1_credit_1_grant,
    input  io_outChannels_1_credit_0_grant,
    output[54:0] io_outChannels_0_flit_x,
    output io_outChannels_0_flitValid,
    input  io_outChannels_0_credit_1_grant,
    input  io_outChannels_0_credit_0_grant,
    output[31:0] io_counters_1_counterVal,
    output[7:0] io_counters_1_counterIndex,
    output[31:0] io_counters_0_counterVal,
    output[7:0] io_counters_0_counterIndex,
    input  io_bypass
);

  wire bp_io_x_inChannels_4_credit_1_grant;
  wire bp_io_x_inChannels_4_credit_0_grant;
  wire bp_io_x_inChannels_3_credit_1_grant;
  wire bp_io_x_inChannels_3_credit_0_grant;
  wire bp_io_x_inChannels_2_credit_1_grant;
  wire bp_io_x_inChannels_2_credit_0_grant;
  wire bp_io_x_inChannels_1_credit_1_grant;
  wire bp_io_x_inChannels_1_credit_0_grant;
  wire bp_io_x_inChannels_0_credit_1_grant;
  wire bp_io_x_inChannels_0_credit_0_grant;
  wire[54:0] bp_io_x_outChannels_4_flit_x;
  wire bp_io_x_outChannels_4_flitValid;
  wire[54:0] bp_io_x_outChannels_3_flit_x;
  wire bp_io_x_outChannels_3_flitValid;
  wire[54:0] bp_io_x_outChannels_2_flit_x;
  wire bp_io_x_outChannels_2_flitValid;
  wire[54:0] bp_io_x_outChannels_1_flit_x;
  wire bp_io_x_outChannels_1_flitValid;
  wire[54:0] bp_io_x_outChannels_0_flit_x;
  wire bp_io_x_outChannels_0_flitValid;
  wire[31:0] bp_io_x_counters_1_counterVal;
  wire[7:0] bp_io_x_counters_1_counterIndex;
  wire[31:0] bp_io_x_counters_0_counterVal;
  wire[7:0] bp_io_x_counters_0_counterIndex;
  wire[54:0] bp_io_y_inChannels_4_flit_x;
  wire bp_io_y_inChannels_4_flitValid;
  wire[54:0] bp_io_y_inChannels_3_flit_x;
  wire bp_io_y_inChannels_3_flitValid;
  wire[54:0] bp_io_y_inChannels_2_flit_x;
  wire bp_io_y_inChannels_2_flitValid;
  wire[54:0] bp_io_y_inChannels_1_flit_x;
  wire bp_io_y_inChannels_1_flitValid;
  wire[54:0] bp_io_y_inChannels_0_flit_x;
  wire bp_io_y_inChannels_0_flitValid;
  wire bp_io_y_outChannels_4_credit_1_grant;
  wire bp_io_y_outChannels_4_credit_0_grant;
  wire bp_io_y_outChannels_3_credit_1_grant;
  wire bp_io_y_outChannels_3_credit_0_grant;
  wire bp_io_y_outChannels_2_credit_1_grant;
  wire bp_io_y_outChannels_2_credit_0_grant;
  wire bp_io_y_outChannels_1_credit_1_grant;
  wire bp_io_y_outChannels_1_credit_0_grant;
  wire bp_io_y_outChannels_0_credit_1_grant;
  wire bp_io_y_outChannels_0_credit_0_grant;
  wire x_io_inChannels_4_credit_1_grant;
  wire x_io_inChannels_4_credit_0_grant;
  wire x_io_inChannels_3_credit_1_grant;
  wire x_io_inChannels_3_credit_0_grant;
  wire x_io_inChannels_2_credit_1_grant;
  wire x_io_inChannels_2_credit_0_grant;
  wire x_io_inChannels_1_credit_1_grant;
  wire x_io_inChannels_1_credit_0_grant;
  wire x_io_inChannels_0_credit_1_grant;
  wire x_io_inChannels_0_credit_0_grant;
  wire[54:0] x_io_outChannels_4_flit_x;
  wire x_io_outChannels_4_flitValid;
  wire[54:0] x_io_outChannels_3_flit_x;
  wire x_io_outChannels_3_flitValid;
  wire[54:0] x_io_outChannels_2_flit_x;
  wire x_io_outChannels_2_flitValid;
  wire[54:0] x_io_outChannels_1_flit_x;
  wire x_io_outChannels_1_flitValid;
  wire[54:0] x_io_outChannels_0_flit_x;
  wire x_io_outChannels_0_flitValid;
  wire[31:0] x_io_counters_0_counterVal;


  assign io_counters_0_counterIndex = bp_io_x_counters_0_counterIndex;
  assign io_counters_0_counterVal = bp_io_x_counters_0_counterVal;
  assign io_counters_1_counterIndex = bp_io_x_counters_1_counterIndex;
  assign io_counters_1_counterVal = bp_io_x_counters_1_counterVal;
  assign io_outChannels_0_flitValid = bp_io_x_outChannels_0_flitValid;
  assign io_outChannels_0_flit_x = bp_io_x_outChannels_0_flit_x;
  assign io_outChannels_1_flitValid = bp_io_x_outChannels_1_flitValid;
  assign io_outChannels_1_flit_x = bp_io_x_outChannels_1_flit_x;
  assign io_outChannels_2_flitValid = bp_io_x_outChannels_2_flitValid;
  assign io_outChannels_2_flit_x = bp_io_x_outChannels_2_flit_x;
  assign io_outChannels_3_flitValid = bp_io_x_outChannels_3_flitValid;
  assign io_outChannels_3_flit_x = bp_io_x_outChannels_3_flit_x;
  assign io_outChannels_4_flitValid = bp_io_x_outChannels_4_flitValid;
  assign io_outChannels_4_flit_x = bp_io_x_outChannels_4_flit_x;
  assign io_inChannels_0_credit_0_grant = bp_io_x_inChannels_0_credit_0_grant;
  assign io_inChannels_0_credit_1_grant = bp_io_x_inChannels_0_credit_1_grant;
  assign io_inChannels_1_credit_0_grant = bp_io_x_inChannels_1_credit_0_grant;
  assign io_inChannels_1_credit_1_grant = bp_io_x_inChannels_1_credit_1_grant;
  assign io_inChannels_2_credit_0_grant = bp_io_x_inChannels_2_credit_0_grant;
  assign io_inChannels_2_credit_1_grant = bp_io_x_inChannels_2_credit_1_grant;
  assign io_inChannels_3_credit_0_grant = bp_io_x_inChannels_3_credit_0_grant;
  assign io_inChannels_3_credit_1_grant = bp_io_x_inChannels_3_credit_1_grant;
  assign io_inChannels_4_credit_0_grant = bp_io_x_inChannels_4_credit_0_grant;
  assign io_inChannels_4_credit_1_grant = bp_io_x_inChannels_4_credit_1_grant;
  wire clkOut;
  VCRouterBypass bp(.clk(clk), .reset(reset),
       .io_x_inChannels_4_flit_x( io_inChannels_4_flit_x ),
       .io_x_inChannels_4_flitValid( io_inChannels_4_flitValid ),
       .io_x_inChannels_4_credit_1_grant( bp_io_x_inChannels_4_credit_1_grant ),
       .io_x_inChannels_4_credit_0_grant( bp_io_x_inChannels_4_credit_0_grant ),
       .io_x_inChannels_3_flit_x( io_inChannels_3_flit_x ),
       .io_x_inChannels_3_flitValid( io_inChannels_3_flitValid ),
       .io_x_inChannels_3_credit_1_grant( bp_io_x_inChannels_3_credit_1_grant ),
       .io_x_inChannels_3_credit_0_grant( bp_io_x_inChannels_3_credit_0_grant ),
       .io_x_inChannels_2_flit_x( io_inChannels_2_flit_x ),
       .io_x_inChannels_2_flitValid( io_inChannels_2_flitValid ),
       .io_x_inChannels_2_credit_1_grant( bp_io_x_inChannels_2_credit_1_grant ),
       .io_x_inChannels_2_credit_0_grant( bp_io_x_inChannels_2_credit_0_grant ),
       .io_x_inChannels_1_flit_x( io_inChannels_1_flit_x ),
       .io_x_inChannels_1_flitValid( io_inChannels_1_flitValid ),
       .io_x_inChannels_1_credit_1_grant( bp_io_x_inChannels_1_credit_1_grant ),
       .io_x_inChannels_1_credit_0_grant( bp_io_x_inChannels_1_credit_0_grant ),
       .io_x_inChannels_0_flit_x( io_inChannels_0_flit_x ),
       .io_x_inChannels_0_flitValid( io_inChannels_0_flitValid ),
       .io_x_inChannels_0_credit_1_grant( bp_io_x_inChannels_0_credit_1_grant ),
       .io_x_inChannels_0_credit_0_grant( bp_io_x_inChannels_0_credit_0_grant ),
       .io_x_outChannels_4_flit_x( bp_io_x_outChannels_4_flit_x ),
       .io_x_outChannels_4_flitValid( bp_io_x_outChannels_4_flitValid ),
       .io_x_outChannels_4_credit_1_grant( io_outChannels_4_credit_1_grant ),
       .io_x_outChannels_4_credit_0_grant( io_outChannels_4_credit_0_grant ),
       .io_x_outChannels_3_flit_x( bp_io_x_outChannels_3_flit_x ),
       .io_x_outChannels_3_flitValid( bp_io_x_outChannels_3_flitValid ),
       .io_x_outChannels_3_credit_1_grant( io_outChannels_3_credit_1_grant ),
       .io_x_outChannels_3_credit_0_grant( io_outChannels_3_credit_0_grant ),
       .io_x_outChannels_2_flit_x( bp_io_x_outChannels_2_flit_x ),
       .io_x_outChannels_2_flitValid( bp_io_x_outChannels_2_flitValid ),
       .io_x_outChannels_2_credit_1_grant( io_outChannels_2_credit_1_grant ),
       .io_x_outChannels_2_credit_0_grant( io_outChannels_2_credit_0_grant ),
       .io_x_outChannels_1_flit_x( bp_io_x_outChannels_1_flit_x ),
       .io_x_outChannels_1_flitValid( bp_io_x_outChannels_1_flitValid ),
       .io_x_outChannels_1_credit_1_grant( io_outChannels_1_credit_1_grant ),
       .io_x_outChannels_1_credit_0_grant( io_outChannels_1_credit_0_grant ),
       .io_x_outChannels_0_flit_x( bp_io_x_outChannels_0_flit_x ),
       .io_x_outChannels_0_flitValid( bp_io_x_outChannels_0_flitValid ),
       .io_x_outChannels_0_credit_1_grant( io_outChannels_0_credit_1_grant ),
       .io_x_outChannels_0_credit_0_grant( io_outChannels_0_credit_0_grant ),
       .io_x_counters_1_counterVal( bp_io_x_counters_1_counterVal ),
       .io_x_counters_1_counterIndex( bp_io_x_counters_1_counterIndex ),
       .io_x_counters_0_counterVal( bp_io_x_counters_0_counterVal ),
       .io_x_counters_0_counterIndex( bp_io_x_counters_0_counterIndex ),
       .io_y_inChannels_4_flit_x( bp_io_y_inChannels_4_flit_x ),
       .io_y_inChannels_4_flitValid( bp_io_y_inChannels_4_flitValid ),
       .io_y_inChannels_4_credit_1_grant( x_io_inChannels_4_credit_1_grant ),
       .io_y_inChannels_4_credit_0_grant( x_io_inChannels_4_credit_0_grant ),
       .io_y_inChannels_3_flit_x( bp_io_y_inChannels_3_flit_x ),
       .io_y_inChannels_3_flitValid( bp_io_y_inChannels_3_flitValid ),
       .io_y_inChannels_3_credit_1_grant( x_io_inChannels_3_credit_1_grant ),
       .io_y_inChannels_3_credit_0_grant( x_io_inChannels_3_credit_0_grant ),
       .io_y_inChannels_2_flit_x( bp_io_y_inChannels_2_flit_x ),
       .io_y_inChannels_2_flitValid( bp_io_y_inChannels_2_flitValid ),
       .io_y_inChannels_2_credit_1_grant( x_io_inChannels_2_credit_1_grant ),
       .io_y_inChannels_2_credit_0_grant( x_io_inChannels_2_credit_0_grant ),
       .io_y_inChannels_1_flit_x( bp_io_y_inChannels_1_flit_x ),
       .io_y_inChannels_1_flitValid( bp_io_y_inChannels_1_flitValid ),
       .io_y_inChannels_1_credit_1_grant( x_io_inChannels_1_credit_1_grant ),
       .io_y_inChannels_1_credit_0_grant( x_io_inChannels_1_credit_0_grant ),
       .io_y_inChannels_0_flit_x( bp_io_y_inChannels_0_flit_x ),
       .io_y_inChannels_0_flitValid( bp_io_y_inChannels_0_flitValid ),
       .io_y_inChannels_0_credit_1_grant( x_io_inChannels_0_credit_1_grant ),
       .io_y_inChannels_0_credit_0_grant( x_io_inChannels_0_credit_0_grant ),
       .io_y_outChannels_4_flit_x( x_io_outChannels_4_flit_x ),
       .io_y_outChannels_4_flitValid( x_io_outChannels_4_flitValid ),
       .io_y_outChannels_4_credit_1_grant( bp_io_y_outChannels_4_credit_1_grant ),
       .io_y_outChannels_4_credit_0_grant( bp_io_y_outChannels_4_credit_0_grant ),
       .io_y_outChannels_3_flit_x( x_io_outChannels_3_flit_x ),
       .io_y_outChannels_3_flitValid( x_io_outChannels_3_flitValid ),
       .io_y_outChannels_3_credit_1_grant( bp_io_y_outChannels_3_credit_1_grant ),
       .io_y_outChannels_3_credit_0_grant( bp_io_y_outChannels_3_credit_0_grant ),
       .io_y_outChannels_2_flit_x( x_io_outChannels_2_flit_x ),
       .io_y_outChannels_2_flitValid( x_io_outChannels_2_flitValid ),
       .io_y_outChannels_2_credit_1_grant( bp_io_y_outChannels_2_credit_1_grant ),
       .io_y_outChannels_2_credit_0_grant( bp_io_y_outChannels_2_credit_0_grant ),
       .io_y_outChannels_1_flit_x( x_io_outChannels_1_flit_x ),
       .io_y_outChannels_1_flitValid( x_io_outChannels_1_flitValid ),
       .io_y_outChannels_1_credit_1_grant( bp_io_y_outChannels_1_credit_1_grant ),
       .io_y_outChannels_1_credit_0_grant( bp_io_y_outChannels_1_credit_0_grant ),
       .io_y_outChannels_0_flit_x( x_io_outChannels_0_flit_x ),
       .io_y_outChannels_0_flitValid( x_io_outChannels_0_flitValid ),
       .io_y_outChannels_0_credit_1_grant( bp_io_y_outChannels_0_credit_1_grant ),
       .io_y_outChannels_0_credit_0_grant( bp_io_y_outChannels_0_credit_0_grant ),
       //.io_y_counters_1_counterVal(  )
       //.io_y_counters_1_counterIndex(  )
       .io_y_counters_0_counterVal( x_io_counters_0_counterVal ),
       //.io_y_counters_0_counterIndex(  )
       .io_bypass( io_bypass ),
       .io_clkOut(clkOut)
  );
  SimpleVCRouter_2 x(.clk(clkOut), .reset(reset),
       .io_inChannels_4_flit_x( bp_io_y_inChannels_4_flit_x ),
       .io_inChannels_4_flitValid( bp_io_y_inChannels_4_flitValid ),
       .io_inChannels_4_credit_1_grant( x_io_inChannels_4_credit_1_grant ),
       .io_inChannels_4_credit_0_grant( x_io_inChannels_4_credit_0_grant ),
       .io_inChannels_3_flit_x( bp_io_y_inChannels_3_flit_x ),
       .io_inChannels_3_flitValid( bp_io_y_inChannels_3_flitValid ),
       .io_inChannels_3_credit_1_grant( x_io_inChannels_3_credit_1_grant ),
       .io_inChannels_3_credit_0_grant( x_io_inChannels_3_credit_0_grant ),
       .io_inChannels_2_flit_x( bp_io_y_inChannels_2_flit_x ),
       .io_inChannels_2_flitValid( bp_io_y_inChannels_2_flitValid ),
       .io_inChannels_2_credit_1_grant( x_io_inChannels_2_credit_1_grant ),
       .io_inChannels_2_credit_0_grant( x_io_inChannels_2_credit_0_grant ),
       .io_inChannels_1_flit_x( bp_io_y_inChannels_1_flit_x ),
       .io_inChannels_1_flitValid( bp_io_y_inChannels_1_flitValid ),
       .io_inChannels_1_credit_1_grant( x_io_inChannels_1_credit_1_grant ),
       .io_inChannels_1_credit_0_grant( x_io_inChannels_1_credit_0_grant ),
       .io_inChannels_0_flit_x( bp_io_y_inChannels_0_flit_x ),
       .io_inChannels_0_flitValid( bp_io_y_inChannels_0_flitValid ),
       .io_inChannels_0_credit_1_grant( x_io_inChannels_0_credit_1_grant ),
       .io_inChannels_0_credit_0_grant( x_io_inChannels_0_credit_0_grant ),
       .io_outChannels_4_flit_x( x_io_outChannels_4_flit_x ),
       .io_outChannels_4_flitValid( x_io_outChannels_4_flitValid ),
       .io_outChannels_4_credit_1_grant( bp_io_y_outChannels_4_credit_1_grant ),
       .io_outChannels_4_credit_0_grant( bp_io_y_outChannels_4_credit_0_grant ),
       .io_outChannels_3_flit_x( x_io_outChannels_3_flit_x ),
       .io_outChannels_3_flitValid( x_io_outChannels_3_flitValid ),
       .io_outChannels_3_credit_1_grant( bp_io_y_outChannels_3_credit_1_grant ),
       .io_outChannels_3_credit_0_grant( bp_io_y_outChannels_3_credit_0_grant ),
       .io_outChannels_2_flit_x( x_io_outChannels_2_flit_x ),
       .io_outChannels_2_flitValid( x_io_outChannels_2_flitValid ),
       .io_outChannels_2_credit_1_grant( bp_io_y_outChannels_2_credit_1_grant ),
       .io_outChannels_2_credit_0_grant( bp_io_y_outChannels_2_credit_0_grant ),
       .io_outChannels_1_flit_x( x_io_outChannels_1_flit_x ),
       .io_outChannels_1_flitValid( x_io_outChannels_1_flitValid ),
       .io_outChannels_1_credit_1_grant( bp_io_y_outChannels_1_credit_1_grant ),
       .io_outChannels_1_credit_0_grant( bp_io_y_outChannels_1_credit_0_grant ),
       .io_outChannels_0_flit_x( x_io_outChannels_0_flit_x ),
       .io_outChannels_0_flitValid( x_io_outChannels_0_flitValid ),
       .io_outChannels_0_credit_1_grant( bp_io_y_outChannels_0_credit_1_grant ),
       .io_outChannels_0_credit_0_grant( bp_io_y_outChannels_0_credit_0_grant ),
       //.io_counters_1_counterVal(  )
       //.io_counters_1_counterIndex(  )
       .io_counters_0_counterVal( x_io_counters_0_counterVal )
       //.io_counters_0_counterIndex(  )
       //.io_bypass(  )
  );
endmodule

module BusProbe_2(input clk, input reset,
    //input [54:0] io_inFlit_4_x
    //input [54:0] io_inFlit_3_x
    input [54:0] io_inFlit_2_x,
    //input [54:0] io_inFlit_1_x
    //input [54:0] io_inFlit_0_x
    input  io_inValid_4,
    input  io_inValid_3,
    input  io_inValid_2,
    input  io_inValid_1,
    input  io_inValid_0,
    input  io_routerCord,
    //input  io_startRecording
    output[15:0] io_cyclesChannelBusy_4,
    output[15:0] io_cyclesChannelBusy_3,
    output[15:0] io_cyclesChannelBusy_2,
    output[15:0] io_cyclesChannelBusy_1,
    output[15:0] io_cyclesChannelBusy_0,
    output[15:0] io_cyclesRouterBusy
);

  reg[0:0] T0;
  reg [15:0] cyclesRouterBusy;
  wire[15:0] T29;
  wire[15:0] T1;
  wire[15:0] T2;
  wire T3;
  wire[4:0] T4;
  wire[4:0] T5;
  wire[2:0] T6;
  wire[1:0] T7;
  reg  cyclesChannelBusyScoreboard_0;
  wire T30;
  wire T8;
  wire T9;
  reg  cyclesChannelBusyScoreboard_1;
  wire T31;
  wire T10;
  wire T11;
  reg  cyclesChannelBusyScoreboard_2;
  wire T32;
  wire T12;
  wire T13;
  wire[1:0] T14;
  reg  cyclesChannelBusyScoreboard_3;
  wire T33;
  wire T15;
  wire T16;
  reg  cyclesChannelBusyScoreboard_4;
  wire T34;
  wire T17;
  wire T18;
  reg [15:0] cyclesChannelBusy_0;
  wire[15:0] T35;
  wire[15:0] T19;
  wire[15:0] T20;
  reg [15:0] cyclesChannelBusy_1;
  wire[15:0] T36;
  wire[15:0] T21;
  wire[15:0] T22;
  reg [15:0] cyclesChannelBusy_2;
  wire[15:0] T37;
  wire[15:0] T23;
  wire[15:0] T24;
  reg [15:0] cyclesChannelBusy_3;
  wire[15:0] T38;
  wire[15:0] T25;
  wire[15:0] T26;
  reg [15:0] cyclesChannelBusy_4;
  wire[15:0] T39;
  wire[15:0] T27;
  wire[15:0] T28;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    T0 = 1'b0;
    cyclesRouterBusy = {1{1'b0}};
    cyclesChannelBusyScoreboard_0 = {1{1'b0}};
    cyclesChannelBusyScoreboard_1 = {1{1'b0}};
    cyclesChannelBusyScoreboard_2 = {1{1'b0}};
    cyclesChannelBusyScoreboard_3 = {1{1'b0}};
    cyclesChannelBusyScoreboard_4 = {1{1'b0}};
    cyclesChannelBusy_0 = {1{1'b0}};
    cyclesChannelBusy_1 = {1{1'b0}};
    cyclesChannelBusy_2 = {1{1'b0}};
    cyclesChannelBusy_3 = {1{1'b0}};
    cyclesChannelBusy_4 = {1{1'b0}};
  end
// synthesis translate_on
`endif

  assign io_cyclesRouterBusy = cyclesRouterBusy;
  assign T29 = reset ? 16'h0 : T1;
  assign T1 = T3 ? T2 : cyclesRouterBusy;
  assign T2 = cyclesRouterBusy + 16'h1;
  assign T3 = T4 != 5'h0;
  assign T4 = T5;
  assign T5 = {T14, T6};
  assign T6 = {cyclesChannelBusyScoreboard_2, T7};
  assign T7 = {cyclesChannelBusyScoreboard_1, cyclesChannelBusyScoreboard_0};
  assign T30 = reset ? 1'h0 : T8;
  assign T8 = T9 == 1'h0;
  assign T9 = io_inValid_0 ^ 1'h1;
  assign T31 = reset ? 1'h0 : T10;
  assign T10 = T11 == 1'h0;
  assign T11 = io_inValid_1 ^ 1'h1;
  assign T32 = reset ? 1'h0 : T12;
  assign T12 = T13 == 1'h0;
  assign T13 = io_inValid_2 ^ 1'h1;
  assign T14 = {cyclesChannelBusyScoreboard_4, cyclesChannelBusyScoreboard_3};
  assign T33 = reset ? 1'h0 : T15;
  assign T15 = T16 == 1'h0;
  assign T16 = io_inValid_3 ^ 1'h1;
  assign T34 = reset ? 1'h0 : T17;
  assign T17 = T18 == 1'h0;
  assign T18 = io_inValid_4 ^ 1'h1;
  assign io_cyclesChannelBusy_0 = cyclesChannelBusy_0;
  assign T35 = reset ? 16'h0 : T19;
  assign T19 = io_inValid_0 ? T20 : cyclesChannelBusy_0;
  assign T20 = cyclesChannelBusy_0 + 16'h1;
  assign io_cyclesChannelBusy_1 = cyclesChannelBusy_1;
  assign T36 = reset ? 16'h0 : T21;
  assign T21 = io_inValid_1 ? T22 : cyclesChannelBusy_1;
  assign T22 = cyclesChannelBusy_1 + 16'h1;
  assign io_cyclesChannelBusy_2 = cyclesChannelBusy_2;
  assign T37 = reset ? 16'h0 : T23;
  assign T23 = io_inValid_2 ? T24 : cyclesChannelBusy_2;
  assign T24 = cyclesChannelBusy_2 + 16'h1;
  assign io_cyclesChannelBusy_3 = cyclesChannelBusy_3;
  assign T38 = reset ? 16'h0 : T25;
  assign T25 = io_inValid_3 ? T26 : cyclesChannelBusy_3;
  assign T26 = cyclesChannelBusy_3 + 16'h1;
  assign io_cyclesChannelBusy_4 = cyclesChannelBusy_4;
  assign T39 = reset ? 16'h0 : T27;
  assign T27 = io_inValid_4 ? T28 : cyclesChannelBusy_4;
  assign T28 = cyclesChannelBusy_4 + 16'h1;

  always @(posedge clk) begin
`ifndef SYNTHESIS
// synthesis translate_off
  if(reset) T0 <= 1'b1;
  if(!1'h1 && T0 && !reset) begin
    $fwrite(32'h80000002, "ASSERTION FAILED: %s\n", "BusProbe: RouterRadix must be > 1");
    $finish;
  end
// synthesis translate_on
`endif
    if(reset) begin
      cyclesRouterBusy <= 16'h0;
    end else if(T3) begin
      cyclesRouterBusy <= T2;
    end
    if(reset) begin
      cyclesChannelBusyScoreboard_0 <= 1'h0;
    end else begin
      cyclesChannelBusyScoreboard_0 <= T8;
    end
    if(reset) begin
      cyclesChannelBusyScoreboard_1 <= 1'h0;
    end else begin
      cyclesChannelBusyScoreboard_1 <= T10;
    end
    if(reset) begin
      cyclesChannelBusyScoreboard_2 <= 1'h0;
    end else begin
      cyclesChannelBusyScoreboard_2 <= T12;
    end
    if(reset) begin
      cyclesChannelBusyScoreboard_3 <= 1'h0;
    end else begin
      cyclesChannelBusyScoreboard_3 <= T15;
    end
    if(reset) begin
      cyclesChannelBusyScoreboard_4 <= 1'h0;
    end else begin
      cyclesChannelBusyScoreboard_4 <= T17;
    end
    if(reset) begin
      cyclesChannelBusy_0 <= 16'h0;
    end else if(io_inValid_0) begin
      cyclesChannelBusy_0 <= T20;
    end
    if(reset) begin
      cyclesChannelBusy_1 <= 16'h0;
    end else if(io_inValid_1) begin
      cyclesChannelBusy_1 <= T22;
    end
    if(reset) begin
      cyclesChannelBusy_2 <= 16'h0;
    end else if(io_inValid_2) begin
      cyclesChannelBusy_2 <= T24;
    end
    if(reset) begin
      cyclesChannelBusy_3 <= 16'h0;
    end else if(io_inValid_3) begin
      cyclesChannelBusy_3 <= T26;
    end
    if(reset) begin
      cyclesChannelBusy_4 <= 16'h0;
    end else if(io_inValid_4) begin
      cyclesChannelBusy_4 <= T28;
    end
  end
endmodule

module OpenSoC_VCConstantEndpoint_0(
    //input [54:0] io_inChannels_4_flit_x
    //input  io_inChannels_4_flitValid
    //output io_inChannels_4_credit_1_grant
    //output io_inChannels_4_credit_0_grant
    //input [54:0] io_inChannels_3_flit_x
    //input  io_inChannels_3_flitValid
    //output io_inChannels_3_credit_1_grant
    //output io_inChannels_3_credit_0_grant
    //input [54:0] io_inChannels_2_flit_x
    //input  io_inChannels_2_flitValid
    //output io_inChannels_2_credit_1_grant
    //output io_inChannels_2_credit_0_grant
    input [54:0] io_inChannels_1_flit_x,
    input  io_inChannels_1_flitValid,
    //output io_inChannels_1_credit_1_grant
    //output io_inChannels_1_credit_0_grant
    //input [54:0] io_inChannels_0_flit_x
    //input  io_inChannels_0_flitValid
    //output io_inChannels_0_credit_1_grant
    //output io_inChannels_0_credit_0_grant
    output[54:0] io_outChannels_4_flit_x,
    output io_outChannels_4_flitValid,
    //input  io_outChannels_4_credit_1_grant
    //input  io_outChannels_4_credit_0_grant
    output[54:0] io_outChannels_3_flit_x,
    output io_outChannels_3_flitValid,
    //input  io_outChannels_3_credit_1_grant
    //input  io_outChannels_3_credit_0_grant
    output[54:0] io_outChannels_2_flit_x,
    output io_outChannels_2_flitValid,
    //input  io_outChannels_2_credit_1_grant
    //input  io_outChannels_2_credit_0_grant
    output[54:0] io_outChannels_1_flit_x,
    output io_outChannels_1_flitValid,
    input  io_outChannels_1_credit_1_grant,
    input  io_outChannels_1_credit_0_grant,
    output[54:0] io_outChannels_0_flit_x,
    output io_outChannels_0_flitValid
    //input  io_outChannels_0_credit_1_grant
    //input  io_outChannels_0_credit_0_grant
    //output[31:0] io_counters_1_counterVal
    //output[7:0] io_counters_1_counterIndex
    //output[31:0] io_counters_0_counterVal
    //output[7:0] io_counters_0_counterIndex
    //input  io_bypass
);

  wire[54:0] T0;
  wire[54:0] T1;
  wire[54:0] T2;
  wire[54:0] T3;
  wire[54:0] T4;


`ifndef SYNTHESIS
// synthesis translate_off
//  assign io_counters_0_counterIndex = {1{1'b0}};
//  assign io_counters_0_counterVal = {1{1'b0}};
//  assign io_counters_1_counterIndex = {1{1'b0}};
//  assign io_counters_1_counterVal = {1{1'b0}};
//  assign io_inChannels_0_credit_0_grant = {1{1'b0}};
//  assign io_inChannels_0_credit_1_grant = {1{1'b0}};
//  assign io_inChannels_1_credit_0_grant = {1{1'b0}};
//  assign io_inChannels_1_credit_1_grant = {1{1'b0}};
//  assign io_inChannels_2_credit_0_grant = {1{1'b0}};
//  assign io_inChannels_2_credit_1_grant = {1{1'b0}};
//  assign io_inChannels_3_credit_0_grant = {1{1'b0}};
//  assign io_inChannels_3_credit_1_grant = {1{1'b0}};
//  assign io_inChannels_4_credit_0_grant = {1{1'b0}};
//  assign io_inChannels_4_credit_1_grant = {1{1'b0}};
// synthesis translate_on
`endif
  assign io_outChannels_0_flitValid = 1'h0;
  assign io_outChannels_0_flit_x = T0;
  assign T0 = 55'h0;
  assign io_outChannels_1_flitValid = 1'h0;
  assign io_outChannels_1_flit_x = T1;
  assign T1 = 55'h0;
  assign io_outChannels_2_flitValid = 1'h0;
  assign io_outChannels_2_flit_x = T2;
  assign T2 = 55'h0;
  assign io_outChannels_3_flitValid = 1'h0;
  assign io_outChannels_3_flit_x = T3;
  assign T3 = 55'h0;
  assign io_outChannels_4_flitValid = 1'h0;
  assign io_outChannels_4_flit_x = T4;
  assign T4 = 55'h0;
endmodule

module OpenSoC_VCConstantEndpoint_1(
    //input [54:0] io_inChannels_4_flit_x
    //input  io_inChannels_4_flitValid
    //output io_inChannels_4_credit_1_grant
    //output io_inChannels_4_credit_0_grant
    input [54:0] io_inChannels_3_flit_x,
    input  io_inChannels_3_flitValid,
    //output io_inChannels_3_credit_1_grant
    //output io_inChannels_3_credit_0_grant
    //input [54:0] io_inChannels_2_flit_x
    //input  io_inChannels_2_flitValid
    //output io_inChannels_2_credit_1_grant
    //output io_inChannels_2_credit_0_grant
    //input [54:0] io_inChannels_1_flit_x
    //input  io_inChannels_1_flitValid
    //output io_inChannels_1_credit_1_grant
    //output io_inChannels_1_credit_0_grant
    //input [54:0] io_inChannels_0_flit_x
    //input  io_inChannels_0_flitValid
    //output io_inChannels_0_credit_1_grant
    //output io_inChannels_0_credit_0_grant
    output[54:0] io_outChannels_4_flit_x,
    output io_outChannels_4_flitValid,
    //input  io_outChannels_4_credit_1_grant
    //input  io_outChannels_4_credit_0_grant
    output[54:0] io_outChannels_3_flit_x,
    output io_outChannels_3_flitValid,
    input  io_outChannels_3_credit_1_grant,
    input  io_outChannels_3_credit_0_grant,
    output[54:0] io_outChannels_2_flit_x,
    output io_outChannels_2_flitValid,
    //input  io_outChannels_2_credit_1_grant
    //input  io_outChannels_2_credit_0_grant
    output[54:0] io_outChannels_1_flit_x,
    output io_outChannels_1_flitValid,
    //input  io_outChannels_1_credit_1_grant
    //input  io_outChannels_1_credit_0_grant
    output[54:0] io_outChannels_0_flit_x,
    output io_outChannels_0_flitValid
    //input  io_outChannels_0_credit_1_grant
    //input  io_outChannels_0_credit_0_grant
    //output[31:0] io_counters_1_counterVal
    //output[7:0] io_counters_1_counterIndex
    //output[31:0] io_counters_0_counterVal
    //output[7:0] io_counters_0_counterIndex
    //input  io_bypass
);

  wire[54:0] T0;
  wire[54:0] T1;
  wire[54:0] T2;
  wire[54:0] T3;
  wire[54:0] T4;


`ifndef SYNTHESIS
// synthesis translate_off
//  assign io_counters_0_counterIndex = {1{1'b0}};
//  assign io_counters_0_counterVal = {1{1'b0}};
//  assign io_counters_1_counterIndex = {1{1'b0}};
//  assign io_counters_1_counterVal = {1{1'b0}};
//  assign io_inChannels_0_credit_0_grant = {1{1'b0}};
//  assign io_inChannels_0_credit_1_grant = {1{1'b0}};
//  assign io_inChannels_1_credit_0_grant = {1{1'b0}};
//  assign io_inChannels_1_credit_1_grant = {1{1'b0}};
//  assign io_inChannels_2_credit_0_grant = {1{1'b0}};
//  assign io_inChannels_2_credit_1_grant = {1{1'b0}};
//  assign io_inChannels_3_credit_0_grant = {1{1'b0}};
//  assign io_inChannels_3_credit_1_grant = {1{1'b0}};
//  assign io_inChannels_4_credit_0_grant = {1{1'b0}};
//  assign io_inChannels_4_credit_1_grant = {1{1'b0}};
// synthesis translate_on
`endif
  assign io_outChannels_0_flitValid = 1'h0;
  assign io_outChannels_0_flit_x = T0;
  assign T0 = 55'h0;
  assign io_outChannels_1_flitValid = 1'h0;
  assign io_outChannels_1_flit_x = T1;
  assign T1 = 55'h0;
  assign io_outChannels_2_flitValid = 1'h0;
  assign io_outChannels_2_flit_x = T2;
  assign T2 = 55'h0;
  assign io_outChannels_3_flitValid = 1'h0;
  assign io_outChannels_3_flit_x = T3;
  assign T3 = 55'h0;
  assign io_outChannels_4_flitValid = 1'h0;
  assign io_outChannels_4_flit_x = T4;
  assign T4 = 55'h0;
endmodule

module OpenSoC_VCConstantEndpoint_2(
    input [54:0] io_inChannels_4_flit_x,
    input  io_inChannels_4_flitValid,
    //output io_inChannels_4_credit_1_grant
    //output io_inChannels_4_credit_0_grant
    //input [54:0] io_inChannels_3_flit_x
    //input  io_inChannels_3_flitValid
    //output io_inChannels_3_credit_1_grant
    //output io_inChannels_3_credit_0_grant
    //input [54:0] io_inChannels_2_flit_x
    //input  io_inChannels_2_flitValid
    //output io_inChannels_2_credit_1_grant
    //output io_inChannels_2_credit_0_grant
    //input [54:0] io_inChannels_1_flit_x
    //input  io_inChannels_1_flitValid
    //output io_inChannels_1_credit_1_grant
    //output io_inChannels_1_credit_0_grant
    //input [54:0] io_inChannels_0_flit_x
    //input  io_inChannels_0_flitValid
    //output io_inChannels_0_credit_1_grant
    //output io_inChannels_0_credit_0_grant
    output[54:0] io_outChannels_4_flit_x,
    output io_outChannels_4_flitValid,
    input  io_outChannels_4_credit_1_grant,
    input  io_outChannels_4_credit_0_grant,
    output[54:0] io_outChannels_3_flit_x,
    output io_outChannels_3_flitValid,
    //input  io_outChannels_3_credit_1_grant
    //input  io_outChannels_3_credit_0_grant
    output[54:0] io_outChannels_2_flit_x,
    output io_outChannels_2_flitValid,
    //input  io_outChannels_2_credit_1_grant
    //input  io_outChannels_2_credit_0_grant
    output[54:0] io_outChannels_1_flit_x,
    output io_outChannels_1_flitValid,
    //input  io_outChannels_1_credit_1_grant
    //input  io_outChannels_1_credit_0_grant
    output[54:0] io_outChannels_0_flit_x,
    output io_outChannels_0_flitValid
    //input  io_outChannels_0_credit_1_grant
    //input  io_outChannels_0_credit_0_grant
    //output[31:0] io_counters_1_counterVal
    //output[7:0] io_counters_1_counterIndex
    //output[31:0] io_counters_0_counterVal
    //output[7:0] io_counters_0_counterIndex
    //input  io_bypass
);

  wire[54:0] T0;
  wire[54:0] T1;
  wire[54:0] T2;
  wire[54:0] T3;
  wire[54:0] T4;


`ifndef SYNTHESIS
// synthesis translate_off
//  assign io_counters_0_counterIndex = {1{1'b0}};
//  assign io_counters_0_counterVal = {1{1'b0}};
//  assign io_counters_1_counterIndex = {1{1'b0}};
//  assign io_counters_1_counterVal = {1{1'b0}};
//  assign io_inChannels_0_credit_0_grant = {1{1'b0}};
//  assign io_inChannels_0_credit_1_grant = {1{1'b0}};
//  assign io_inChannels_1_credit_0_grant = {1{1'b0}};
//  assign io_inChannels_1_credit_1_grant = {1{1'b0}};
//  assign io_inChannels_2_credit_0_grant = {1{1'b0}};
//  assign io_inChannels_2_credit_1_grant = {1{1'b0}};
//  assign io_inChannels_3_credit_0_grant = {1{1'b0}};
//  assign io_inChannels_3_credit_1_grant = {1{1'b0}};
//  assign io_inChannels_4_credit_0_grant = {1{1'b0}};
//  assign io_inChannels_4_credit_1_grant = {1{1'b0}};
// synthesis translate_on
`endif
  assign io_outChannels_0_flitValid = 1'h0;
  assign io_outChannels_0_flit_x = T0;
  assign T0 = 55'h0;
  assign io_outChannels_1_flitValid = 1'h0;
  assign io_outChannels_1_flit_x = T1;
  assign T1 = 55'h0;
  assign io_outChannels_2_flitValid = 1'h0;
  assign io_outChannels_2_flit_x = T2;
  assign T2 = 55'h0;
  assign io_outChannels_3_flitValid = 1'h0;
  assign io_outChannels_3_flit_x = T3;
  assign T3 = 55'h0;
  assign io_outChannels_4_flitValid = 1'h0;
  assign io_outChannels_4_flit_x = T4;
  assign T4 = 55'h0;
endmodule

module OpenSoC_VCConstantEndpoint_3(
    //input [54:0] io_inChannels_4_flit_x
    //input  io_inChannels_4_flitValid
    //output io_inChannels_4_credit_1_grant
    //output io_inChannels_4_credit_0_grant
    //input [54:0] io_inChannels_3_flit_x
    //input  io_inChannels_3_flitValid
    //output io_inChannels_3_credit_1_grant
    //output io_inChannels_3_credit_0_grant
    input [54:0] io_inChannels_2_flit_x,
    input  io_inChannels_2_flitValid,
    //output io_inChannels_2_credit_1_grant
    //output io_inChannels_2_credit_0_grant
    //input [54:0] io_inChannels_1_flit_x
    //input  io_inChannels_1_flitValid
    //output io_inChannels_1_credit_1_grant
    //output io_inChannels_1_credit_0_grant
    //input [54:0] io_inChannels_0_flit_x
    //input  io_inChannels_0_flitValid
    //output io_inChannels_0_credit_1_grant
    //output io_inChannels_0_credit_0_grant
    output[54:0] io_outChannels_4_flit_x,
    output io_outChannels_4_flitValid,
    //input  io_outChannels_4_credit_1_grant
    //input  io_outChannels_4_credit_0_grant
    output[54:0] io_outChannels_3_flit_x,
    output io_outChannels_3_flitValid,
    //input  io_outChannels_3_credit_1_grant
    //input  io_outChannels_3_credit_0_grant
    output[54:0] io_outChannels_2_flit_x,
    output io_outChannels_2_flitValid,
    input  io_outChannels_2_credit_1_grant,
    input  io_outChannels_2_credit_0_grant,
    output[54:0] io_outChannels_1_flit_x,
    output io_outChannels_1_flitValid,
    //input  io_outChannels_1_credit_1_grant
    //input  io_outChannels_1_credit_0_grant
    output[54:0] io_outChannels_0_flit_x,
    output io_outChannels_0_flitValid
    //input  io_outChannels_0_credit_1_grant
    //input  io_outChannels_0_credit_0_grant
    //output[31:0] io_counters_1_counterVal
    //output[7:0] io_counters_1_counterIndex
    //output[31:0] io_counters_0_counterVal
    //output[7:0] io_counters_0_counterIndex
    //input  io_bypass
);

  wire[54:0] T0;
  wire[54:0] T1;
  wire[54:0] T2;
  wire[54:0] T3;
  wire[54:0] T4;


`ifndef SYNTHESIS
// synthesis translate_off
//  assign io_counters_0_counterIndex = {1{1'b0}};
//  assign io_counters_0_counterVal = {1{1'b0}};
//  assign io_counters_1_counterIndex = {1{1'b0}};
//  assign io_counters_1_counterVal = {1{1'b0}};
//  assign io_inChannels_0_credit_0_grant = {1{1'b0}};
//  assign io_inChannels_0_credit_1_grant = {1{1'b0}};
//  assign io_inChannels_1_credit_0_grant = {1{1'b0}};
//  assign io_inChannels_1_credit_1_grant = {1{1'b0}};
//  assign io_inChannels_2_credit_0_grant = {1{1'b0}};
//  assign io_inChannels_2_credit_1_grant = {1{1'b0}};
//  assign io_inChannels_3_credit_0_grant = {1{1'b0}};
//  assign io_inChannels_3_credit_1_grant = {1{1'b0}};
//  assign io_inChannels_4_credit_0_grant = {1{1'b0}};
//  assign io_inChannels_4_credit_1_grant = {1{1'b0}};
// synthesis translate_on
`endif
  assign io_outChannels_0_flitValid = 1'h0;
  assign io_outChannels_0_flit_x = T0;
  assign T0 = 55'h0;
  assign io_outChannels_1_flitValid = 1'h0;
  assign io_outChannels_1_flit_x = T1;
  assign T1 = 55'h0;
  assign io_outChannels_2_flitValid = 1'h0;
  assign io_outChannels_2_flit_x = T2;
  assign T2 = 55'h0;
  assign io_outChannels_3_flitValid = 1'h0;
  assign io_outChannels_3_flit_x = T3;
  assign T3 = 55'h0;
  assign io_outChannels_4_flitValid = 1'h0;
  assign io_outChannels_4_flit_x = T4;
  assign T4 = 55'h0;
endmodule

module VCCMesh(input clk, input reset,
    input [54:0] io_inChannels_2_flit_x,
    input  io_inChannels_2_flitValid,
    output io_inChannels_2_credit_1_grant,
    output io_inChannels_2_credit_0_grant,
    input [54:0] io_inChannels_1_flit_x,
    input  io_inChannels_1_flitValid,
    output io_inChannels_1_credit_1_grant,
    output io_inChannels_1_credit_0_grant,
    input [54:0] io_inChannels_0_flit_x,
    input  io_inChannels_0_flitValid,
    output io_inChannels_0_credit_1_grant,
    output io_inChannels_0_credit_0_grant,
    output[54:0] io_outChannels_2_flit_x,
    output io_outChannels_2_flitValid,
    input  io_outChannels_2_credit_1_grant,
    input  io_outChannels_2_credit_0_grant,
    output[54:0] io_outChannels_1_flit_x,
    output io_outChannels_1_flitValid,
    input  io_outChannels_1_credit_1_grant,
    input  io_outChannels_1_credit_0_grant,
    output[54:0] io_outChannels_0_flit_x,
    output io_outChannels_0_flitValid,
    input  io_outChannels_0_credit_1_grant,
    input  io_outChannels_0_credit_0_grant,
    //output[15:0] io_cyclesRouterBusy_127
    //output[15:0] io_cyclesRouterBusy_126
    //output[15:0] io_cyclesRouterBusy_125
    //output[15:0] io_cyclesRouterBusy_124
    //output[15:0] io_cyclesRouterBusy_123
    //output[15:0] io_cyclesRouterBusy_122
    //output[15:0] io_cyclesRouterBusy_121
    //output[15:0] io_cyclesRouterBusy_120
    //output[15:0] io_cyclesRouterBusy_119
    //output[15:0] io_cyclesRouterBusy_118
    //output[15:0] io_cyclesRouterBusy_117
    //output[15:0] io_cyclesRouterBusy_116
    //output[15:0] io_cyclesRouterBusy_115
    //output[15:0] io_cyclesRouterBusy_114
    //output[15:0] io_cyclesRouterBusy_113
    //output[15:0] io_cyclesRouterBusy_112
    //output[15:0] io_cyclesRouterBusy_111
    //output[15:0] io_cyclesRouterBusy_110
    //output[15:0] io_cyclesRouterBusy_109
    //output[15:0] io_cyclesRouterBusy_108
    //output[15:0] io_cyclesRouterBusy_107
    //output[15:0] io_cyclesRouterBusy_106
    //output[15:0] io_cyclesRouterBusy_105
    //output[15:0] io_cyclesRouterBusy_104
    //output[15:0] io_cyclesRouterBusy_103
    //output[15:0] io_cyclesRouterBusy_102
    //output[15:0] io_cyclesRouterBusy_101
    //output[15:0] io_cyclesRouterBusy_100
    //output[15:0] io_cyclesRouterBusy_99
    //output[15:0] io_cyclesRouterBusy_98
    //output[15:0] io_cyclesRouterBusy_97
    //output[15:0] io_cyclesRouterBusy_96
    //output[15:0] io_cyclesRouterBusy_95
    //output[15:0] io_cyclesRouterBusy_94
    //output[15:0] io_cyclesRouterBusy_93
    //output[15:0] io_cyclesRouterBusy_92
    //output[15:0] io_cyclesRouterBusy_91
    //output[15:0] io_cyclesRouterBusy_90
    //output[15:0] io_cyclesRouterBusy_89
    //output[15:0] io_cyclesRouterBusy_88
    //output[15:0] io_cyclesRouterBusy_87
    //output[15:0] io_cyclesRouterBusy_86
    //output[15:0] io_cyclesRouterBusy_85
    //output[15:0] io_cyclesRouterBusy_84
    //output[15:0] io_cyclesRouterBusy_83
    //output[15:0] io_cyclesRouterBusy_82
    //output[15:0] io_cyclesRouterBusy_81
    //output[15:0] io_cyclesRouterBusy_80
    //output[15:0] io_cyclesRouterBusy_79
    //output[15:0] io_cyclesRouterBusy_78
    //output[15:0] io_cyclesRouterBusy_77
    //output[15:0] io_cyclesRouterBusy_76
    //output[15:0] io_cyclesRouterBusy_75
    //output[15:0] io_cyclesRouterBusy_74
    //output[15:0] io_cyclesRouterBusy_73
    //output[15:0] io_cyclesRouterBusy_72
    //output[15:0] io_cyclesRouterBusy_71
    //output[15:0] io_cyclesRouterBusy_70
    //output[15:0] io_cyclesRouterBusy_69
    //output[15:0] io_cyclesRouterBusy_68
    //output[15:0] io_cyclesRouterBusy_67
    //output[15:0] io_cyclesRouterBusy_66
    //output[15:0] io_cyclesRouterBusy_65
    //output[15:0] io_cyclesRouterBusy_64
    //output[15:0] io_cyclesRouterBusy_63
    //output[15:0] io_cyclesRouterBusy_62
    //output[15:0] io_cyclesRouterBusy_61
    //output[15:0] io_cyclesRouterBusy_60
    //output[15:0] io_cyclesRouterBusy_59
    //output[15:0] io_cyclesRouterBusy_58
    //output[15:0] io_cyclesRouterBusy_57
    //output[15:0] io_cyclesRouterBusy_56
    //output[15:0] io_cyclesRouterBusy_55
    //output[15:0] io_cyclesRouterBusy_54
    //output[15:0] io_cyclesRouterBusy_53
    //output[15:0] io_cyclesRouterBusy_52
    //output[15:0] io_cyclesRouterBusy_51
    //output[15:0] io_cyclesRouterBusy_50
    //output[15:0] io_cyclesRouterBusy_49
    //output[15:0] io_cyclesRouterBusy_48
    //output[15:0] io_cyclesRouterBusy_47
    //output[15:0] io_cyclesRouterBusy_46
    //output[15:0] io_cyclesRouterBusy_45
    //output[15:0] io_cyclesRouterBusy_44
    //output[15:0] io_cyclesRouterBusy_43
    //output[15:0] io_cyclesRouterBusy_42
    //output[15:0] io_cyclesRouterBusy_41
    //output[15:0] io_cyclesRouterBusy_40
    //output[15:0] io_cyclesRouterBusy_39
    //output[15:0] io_cyclesRouterBusy_38
    //output[15:0] io_cyclesRouterBusy_37
    //output[15:0] io_cyclesRouterBusy_36
    //output[15:0] io_cyclesRouterBusy_35
    //output[15:0] io_cyclesRouterBusy_34
    //output[15:0] io_cyclesRouterBusy_33
    //output[15:0] io_cyclesRouterBusy_32
    //output[15:0] io_cyclesRouterBusy_31
    //output[15:0] io_cyclesRouterBusy_30
    //output[15:0] io_cyclesRouterBusy_29
    //output[15:0] io_cyclesRouterBusy_28
    //output[15:0] io_cyclesRouterBusy_27
    //output[15:0] io_cyclesRouterBusy_26
    //output[15:0] io_cyclesRouterBusy_25
    //output[15:0] io_cyclesRouterBusy_24
    //output[15:0] io_cyclesRouterBusy_23
    //output[15:0] io_cyclesRouterBusy_22
    //output[15:0] io_cyclesRouterBusy_21
    //output[15:0] io_cyclesRouterBusy_20
    //output[15:0] io_cyclesRouterBusy_19
    //output[15:0] io_cyclesRouterBusy_18
    //output[15:0] io_cyclesRouterBusy_17
    //output[15:0] io_cyclesRouterBusy_16
    //output[15:0] io_cyclesRouterBusy_15
    //output[15:0] io_cyclesRouterBusy_14
    //output[15:0] io_cyclesRouterBusy_13
    //output[15:0] io_cyclesRouterBusy_12
    //output[15:0] io_cyclesRouterBusy_11
    //output[15:0] io_cyclesRouterBusy_10
    //output[15:0] io_cyclesRouterBusy_9
    //output[15:0] io_cyclesRouterBusy_8
    //output[15:0] io_cyclesRouterBusy_7
    //output[15:0] io_cyclesRouterBusy_6
    //output[15:0] io_cyclesRouterBusy_5
    //output[15:0] io_cyclesRouterBusy_4
    //output[15:0] io_cyclesRouterBusy_3
    output[15:0] io_cyclesRouterBusy_2,
    output[15:0] io_cyclesRouterBusy_1,
    output[15:0] io_cyclesRouterBusy_0,
    //output[15:0] io_cyclesChannelBusy_639
    //output[15:0] io_cyclesChannelBusy_638
    //output[15:0] io_cyclesChannelBusy_637
    //output[15:0] io_cyclesChannelBusy_636
    //output[15:0] io_cyclesChannelBusy_635
    //output[15:0] io_cyclesChannelBusy_634
    //output[15:0] io_cyclesChannelBusy_633
    //output[15:0] io_cyclesChannelBusy_632
    //output[15:0] io_cyclesChannelBusy_631
    //output[15:0] io_cyclesChannelBusy_630
    //output[15:0] io_cyclesChannelBusy_629
    //output[15:0] io_cyclesChannelBusy_628
    //output[15:0] io_cyclesChannelBusy_627
    //output[15:0] io_cyclesChannelBusy_626
    //output[15:0] io_cyclesChannelBusy_625
    //output[15:0] io_cyclesChannelBusy_624
    //output[15:0] io_cyclesChannelBusy_623
    //output[15:0] io_cyclesChannelBusy_622
    //output[15:0] io_cyclesChannelBusy_621
    //output[15:0] io_cyclesChannelBusy_620
    //output[15:0] io_cyclesChannelBusy_619
    //output[15:0] io_cyclesChannelBusy_618
    //output[15:0] io_cyclesChannelBusy_617
    //output[15:0] io_cyclesChannelBusy_616
    //output[15:0] io_cyclesChannelBusy_615
    //output[15:0] io_cyclesChannelBusy_614
    //output[15:0] io_cyclesChannelBusy_613
    //output[15:0] io_cyclesChannelBusy_612
    //output[15:0] io_cyclesChannelBusy_611
    //output[15:0] io_cyclesChannelBusy_610
    //output[15:0] io_cyclesChannelBusy_609
    //output[15:0] io_cyclesChannelBusy_608
    //output[15:0] io_cyclesChannelBusy_607
    //output[15:0] io_cyclesChannelBusy_606
    //output[15:0] io_cyclesChannelBusy_605
    //output[15:0] io_cyclesChannelBusy_604
    //output[15:0] io_cyclesChannelBusy_603
    //output[15:0] io_cyclesChannelBusy_602
    //output[15:0] io_cyclesChannelBusy_601
    //output[15:0] io_cyclesChannelBusy_600
    //output[15:0] io_cyclesChannelBusy_599
    //output[15:0] io_cyclesChannelBusy_598
    //output[15:0] io_cyclesChannelBusy_597
    //output[15:0] io_cyclesChannelBusy_596
    //output[15:0] io_cyclesChannelBusy_595
    //output[15:0] io_cyclesChannelBusy_594
    //output[15:0] io_cyclesChannelBusy_593
    //output[15:0] io_cyclesChannelBusy_592
    //output[15:0] io_cyclesChannelBusy_591
    //output[15:0] io_cyclesChannelBusy_590
    //output[15:0] io_cyclesChannelBusy_589
    //output[15:0] io_cyclesChannelBusy_588
    //output[15:0] io_cyclesChannelBusy_587
    //output[15:0] io_cyclesChannelBusy_586
    //output[15:0] io_cyclesChannelBusy_585
    //output[15:0] io_cyclesChannelBusy_584
    //output[15:0] io_cyclesChannelBusy_583
    //output[15:0] io_cyclesChannelBusy_582
    //output[15:0] io_cyclesChannelBusy_581
    //output[15:0] io_cyclesChannelBusy_580
    //output[15:0] io_cyclesChannelBusy_579
    //output[15:0] io_cyclesChannelBusy_578
    //output[15:0] io_cyclesChannelBusy_577
    //output[15:0] io_cyclesChannelBusy_576
    //output[15:0] io_cyclesChannelBusy_575
    //output[15:0] io_cyclesChannelBusy_574
    //output[15:0] io_cyclesChannelBusy_573
    //output[15:0] io_cyclesChannelBusy_572
    //output[15:0] io_cyclesChannelBusy_571
    //output[15:0] io_cyclesChannelBusy_570
    //output[15:0] io_cyclesChannelBusy_569
    //output[15:0] io_cyclesChannelBusy_568
    //output[15:0] io_cyclesChannelBusy_567
    //output[15:0] io_cyclesChannelBusy_566
    //output[15:0] io_cyclesChannelBusy_565
    //output[15:0] io_cyclesChannelBusy_564
    //output[15:0] io_cyclesChannelBusy_563
    //output[15:0] io_cyclesChannelBusy_562
    //output[15:0] io_cyclesChannelBusy_561
    //output[15:0] io_cyclesChannelBusy_560
    //output[15:0] io_cyclesChannelBusy_559
    //output[15:0] io_cyclesChannelBusy_558
    //output[15:0] io_cyclesChannelBusy_557
    //output[15:0] io_cyclesChannelBusy_556
    //output[15:0] io_cyclesChannelBusy_555
    //output[15:0] io_cyclesChannelBusy_554
    //output[15:0] io_cyclesChannelBusy_553
    //output[15:0] io_cyclesChannelBusy_552
    //output[15:0] io_cyclesChannelBusy_551
    //output[15:0] io_cyclesChannelBusy_550
    //output[15:0] io_cyclesChannelBusy_549
    //output[15:0] io_cyclesChannelBusy_548
    //output[15:0] io_cyclesChannelBusy_547
    //output[15:0] io_cyclesChannelBusy_546
    //output[15:0] io_cyclesChannelBusy_545
    //output[15:0] io_cyclesChannelBusy_544
    //output[15:0] io_cyclesChannelBusy_543
    //output[15:0] io_cyclesChannelBusy_542
    //output[15:0] io_cyclesChannelBusy_541
    //output[15:0] io_cyclesChannelBusy_540
    //output[15:0] io_cyclesChannelBusy_539
    //output[15:0] io_cyclesChannelBusy_538
    //output[15:0] io_cyclesChannelBusy_537
    //output[15:0] io_cyclesChannelBusy_536
    //output[15:0] io_cyclesChannelBusy_535
    //output[15:0] io_cyclesChannelBusy_534
    //output[15:0] io_cyclesChannelBusy_533
    //output[15:0] io_cyclesChannelBusy_532
    //output[15:0] io_cyclesChannelBusy_531
    //output[15:0] io_cyclesChannelBusy_530
    //output[15:0] io_cyclesChannelBusy_529
    //output[15:0] io_cyclesChannelBusy_528
    //output[15:0] io_cyclesChannelBusy_527
    //output[15:0] io_cyclesChannelBusy_526
    //output[15:0] io_cyclesChannelBusy_525
    //output[15:0] io_cyclesChannelBusy_524
    //output[15:0] io_cyclesChannelBusy_523
    //output[15:0] io_cyclesChannelBusy_522
    //output[15:0] io_cyclesChannelBusy_521
    //output[15:0] io_cyclesChannelBusy_520
    //output[15:0] io_cyclesChannelBusy_519
    //output[15:0] io_cyclesChannelBusy_518
    //output[15:0] io_cyclesChannelBusy_517
    //output[15:0] io_cyclesChannelBusy_516
    //output[15:0] io_cyclesChannelBusy_515
    //output[15:0] io_cyclesChannelBusy_514
    //output[15:0] io_cyclesChannelBusy_513
    //output[15:0] io_cyclesChannelBusy_512
    //output[15:0] io_cyclesChannelBusy_511
    //output[15:0] io_cyclesChannelBusy_510
    //output[15:0] io_cyclesChannelBusy_509
    //output[15:0] io_cyclesChannelBusy_508
    //output[15:0] io_cyclesChannelBusy_507
    //output[15:0] io_cyclesChannelBusy_506
    //output[15:0] io_cyclesChannelBusy_505
    //output[15:0] io_cyclesChannelBusy_504
    //output[15:0] io_cyclesChannelBusy_503
    //output[15:0] io_cyclesChannelBusy_502
    //output[15:0] io_cyclesChannelBusy_501
    //output[15:0] io_cyclesChannelBusy_500
    //output[15:0] io_cyclesChannelBusy_499
    //output[15:0] io_cyclesChannelBusy_498
    //output[15:0] io_cyclesChannelBusy_497
    //output[15:0] io_cyclesChannelBusy_496
    //output[15:0] io_cyclesChannelBusy_495
    //output[15:0] io_cyclesChannelBusy_494
    //output[15:0] io_cyclesChannelBusy_493
    //output[15:0] io_cyclesChannelBusy_492
    //output[15:0] io_cyclesChannelBusy_491
    //output[15:0] io_cyclesChannelBusy_490
    //output[15:0] io_cyclesChannelBusy_489
    //output[15:0] io_cyclesChannelBusy_488
    //output[15:0] io_cyclesChannelBusy_487
    //output[15:0] io_cyclesChannelBusy_486
    //output[15:0] io_cyclesChannelBusy_485
    //output[15:0] io_cyclesChannelBusy_484
    //output[15:0] io_cyclesChannelBusy_483
    //output[15:0] io_cyclesChannelBusy_482
    //output[15:0] io_cyclesChannelBusy_481
    //output[15:0] io_cyclesChannelBusy_480
    //output[15:0] io_cyclesChannelBusy_479
    //output[15:0] io_cyclesChannelBusy_478
    //output[15:0] io_cyclesChannelBusy_477
    //output[15:0] io_cyclesChannelBusy_476
    //output[15:0] io_cyclesChannelBusy_475
    //output[15:0] io_cyclesChannelBusy_474
    //output[15:0] io_cyclesChannelBusy_473
    //output[15:0] io_cyclesChannelBusy_472
    //output[15:0] io_cyclesChannelBusy_471
    //output[15:0] io_cyclesChannelBusy_470
    //output[15:0] io_cyclesChannelBusy_469
    //output[15:0] io_cyclesChannelBusy_468
    //output[15:0] io_cyclesChannelBusy_467
    //output[15:0] io_cyclesChannelBusy_466
    //output[15:0] io_cyclesChannelBusy_465
    //output[15:0] io_cyclesChannelBusy_464
    //output[15:0] io_cyclesChannelBusy_463
    //output[15:0] io_cyclesChannelBusy_462
    //output[15:0] io_cyclesChannelBusy_461
    //output[15:0] io_cyclesChannelBusy_460
    //output[15:0] io_cyclesChannelBusy_459
    //output[15:0] io_cyclesChannelBusy_458
    //output[15:0] io_cyclesChannelBusy_457
    //output[15:0] io_cyclesChannelBusy_456
    //output[15:0] io_cyclesChannelBusy_455
    //output[15:0] io_cyclesChannelBusy_454
    //output[15:0] io_cyclesChannelBusy_453
    //output[15:0] io_cyclesChannelBusy_452
    //output[15:0] io_cyclesChannelBusy_451
    //output[15:0] io_cyclesChannelBusy_450
    //output[15:0] io_cyclesChannelBusy_449
    //output[15:0] io_cyclesChannelBusy_448
    //output[15:0] io_cyclesChannelBusy_447
    //output[15:0] io_cyclesChannelBusy_446
    //output[15:0] io_cyclesChannelBusy_445
    //output[15:0] io_cyclesChannelBusy_444
    //output[15:0] io_cyclesChannelBusy_443
    //output[15:0] io_cyclesChannelBusy_442
    //output[15:0] io_cyclesChannelBusy_441
    //output[15:0] io_cyclesChannelBusy_440
    //output[15:0] io_cyclesChannelBusy_439
    //output[15:0] io_cyclesChannelBusy_438
    //output[15:0] io_cyclesChannelBusy_437
    //output[15:0] io_cyclesChannelBusy_436
    //output[15:0] io_cyclesChannelBusy_435
    //output[15:0] io_cyclesChannelBusy_434
    //output[15:0] io_cyclesChannelBusy_433
    //output[15:0] io_cyclesChannelBusy_432
    //output[15:0] io_cyclesChannelBusy_431
    //output[15:0] io_cyclesChannelBusy_430
    //output[15:0] io_cyclesChannelBusy_429
    //output[15:0] io_cyclesChannelBusy_428
    //output[15:0] io_cyclesChannelBusy_427
    //output[15:0] io_cyclesChannelBusy_426
    //output[15:0] io_cyclesChannelBusy_425
    //output[15:0] io_cyclesChannelBusy_424
    //output[15:0] io_cyclesChannelBusy_423
    //output[15:0] io_cyclesChannelBusy_422
    //output[15:0] io_cyclesChannelBusy_421
    //output[15:0] io_cyclesChannelBusy_420
    //output[15:0] io_cyclesChannelBusy_419
    //output[15:0] io_cyclesChannelBusy_418
    //output[15:0] io_cyclesChannelBusy_417
    //output[15:0] io_cyclesChannelBusy_416
    //output[15:0] io_cyclesChannelBusy_415
    //output[15:0] io_cyclesChannelBusy_414
    //output[15:0] io_cyclesChannelBusy_413
    //output[15:0] io_cyclesChannelBusy_412
    //output[15:0] io_cyclesChannelBusy_411
    //output[15:0] io_cyclesChannelBusy_410
    //output[15:0] io_cyclesChannelBusy_409
    //output[15:0] io_cyclesChannelBusy_408
    //output[15:0] io_cyclesChannelBusy_407
    //output[15:0] io_cyclesChannelBusy_406
    //output[15:0] io_cyclesChannelBusy_405
    //output[15:0] io_cyclesChannelBusy_404
    //output[15:0] io_cyclesChannelBusy_403
    //output[15:0] io_cyclesChannelBusy_402
    //output[15:0] io_cyclesChannelBusy_401
    //output[15:0] io_cyclesChannelBusy_400
    //output[15:0] io_cyclesChannelBusy_399
    //output[15:0] io_cyclesChannelBusy_398
    //output[15:0] io_cyclesChannelBusy_397
    //output[15:0] io_cyclesChannelBusy_396
    //output[15:0] io_cyclesChannelBusy_395
    //output[15:0] io_cyclesChannelBusy_394
    //output[15:0] io_cyclesChannelBusy_393
    //output[15:0] io_cyclesChannelBusy_392
    //output[15:0] io_cyclesChannelBusy_391
    //output[15:0] io_cyclesChannelBusy_390
    //output[15:0] io_cyclesChannelBusy_389
    //output[15:0] io_cyclesChannelBusy_388
    //output[15:0] io_cyclesChannelBusy_387
    //output[15:0] io_cyclesChannelBusy_386
    //output[15:0] io_cyclesChannelBusy_385
    //output[15:0] io_cyclesChannelBusy_384
    //output[15:0] io_cyclesChannelBusy_383
    //output[15:0] io_cyclesChannelBusy_382
    //output[15:0] io_cyclesChannelBusy_381
    //output[15:0] io_cyclesChannelBusy_380
    //output[15:0] io_cyclesChannelBusy_379
    //output[15:0] io_cyclesChannelBusy_378
    //output[15:0] io_cyclesChannelBusy_377
    //output[15:0] io_cyclesChannelBusy_376
    //output[15:0] io_cyclesChannelBusy_375
    //output[15:0] io_cyclesChannelBusy_374
    //output[15:0] io_cyclesChannelBusy_373
    //output[15:0] io_cyclesChannelBusy_372
    //output[15:0] io_cyclesChannelBusy_371
    //output[15:0] io_cyclesChannelBusy_370
    //output[15:0] io_cyclesChannelBusy_369
    //output[15:0] io_cyclesChannelBusy_368
    //output[15:0] io_cyclesChannelBusy_367
    //output[15:0] io_cyclesChannelBusy_366
    //output[15:0] io_cyclesChannelBusy_365
    //output[15:0] io_cyclesChannelBusy_364
    //output[15:0] io_cyclesChannelBusy_363
    //output[15:0] io_cyclesChannelBusy_362
    //output[15:0] io_cyclesChannelBusy_361
    //output[15:0] io_cyclesChannelBusy_360
    //output[15:0] io_cyclesChannelBusy_359
    //output[15:0] io_cyclesChannelBusy_358
    //output[15:0] io_cyclesChannelBusy_357
    //output[15:0] io_cyclesChannelBusy_356
    //output[15:0] io_cyclesChannelBusy_355
    //output[15:0] io_cyclesChannelBusy_354
    //output[15:0] io_cyclesChannelBusy_353
    //output[15:0] io_cyclesChannelBusy_352
    //output[15:0] io_cyclesChannelBusy_351
    //output[15:0] io_cyclesChannelBusy_350
    //output[15:0] io_cyclesChannelBusy_349
    //output[15:0] io_cyclesChannelBusy_348
    //output[15:0] io_cyclesChannelBusy_347
    //output[15:0] io_cyclesChannelBusy_346
    //output[15:0] io_cyclesChannelBusy_345
    //output[15:0] io_cyclesChannelBusy_344
    //output[15:0] io_cyclesChannelBusy_343
    //output[15:0] io_cyclesChannelBusy_342
    //output[15:0] io_cyclesChannelBusy_341
    //output[15:0] io_cyclesChannelBusy_340
    //output[15:0] io_cyclesChannelBusy_339
    //output[15:0] io_cyclesChannelBusy_338
    //output[15:0] io_cyclesChannelBusy_337
    //output[15:0] io_cyclesChannelBusy_336
    //output[15:0] io_cyclesChannelBusy_335
    //output[15:0] io_cyclesChannelBusy_334
    //output[15:0] io_cyclesChannelBusy_333
    //output[15:0] io_cyclesChannelBusy_332
    //output[15:0] io_cyclesChannelBusy_331
    //output[15:0] io_cyclesChannelBusy_330
    //output[15:0] io_cyclesChannelBusy_329
    //output[15:0] io_cyclesChannelBusy_328
    //output[15:0] io_cyclesChannelBusy_327
    //output[15:0] io_cyclesChannelBusy_326
    //output[15:0] io_cyclesChannelBusy_325
    //output[15:0] io_cyclesChannelBusy_324
    //output[15:0] io_cyclesChannelBusy_323
    //output[15:0] io_cyclesChannelBusy_322
    //output[15:0] io_cyclesChannelBusy_321
    //output[15:0] io_cyclesChannelBusy_320
    //output[15:0] io_cyclesChannelBusy_319
    //output[15:0] io_cyclesChannelBusy_318
    //output[15:0] io_cyclesChannelBusy_317
    //output[15:0] io_cyclesChannelBusy_316
    //output[15:0] io_cyclesChannelBusy_315
    //output[15:0] io_cyclesChannelBusy_314
    //output[15:0] io_cyclesChannelBusy_313
    //output[15:0] io_cyclesChannelBusy_312
    //output[15:0] io_cyclesChannelBusy_311
    //output[15:0] io_cyclesChannelBusy_310
    //output[15:0] io_cyclesChannelBusy_309
    //output[15:0] io_cyclesChannelBusy_308
    //output[15:0] io_cyclesChannelBusy_307
    //output[15:0] io_cyclesChannelBusy_306
    //output[15:0] io_cyclesChannelBusy_305
    //output[15:0] io_cyclesChannelBusy_304
    //output[15:0] io_cyclesChannelBusy_303
    //output[15:0] io_cyclesChannelBusy_302
    //output[15:0] io_cyclesChannelBusy_301
    //output[15:0] io_cyclesChannelBusy_300
    //output[15:0] io_cyclesChannelBusy_299
    //output[15:0] io_cyclesChannelBusy_298
    //output[15:0] io_cyclesChannelBusy_297
    //output[15:0] io_cyclesChannelBusy_296
    //output[15:0] io_cyclesChannelBusy_295
    //output[15:0] io_cyclesChannelBusy_294
    //output[15:0] io_cyclesChannelBusy_293
    //output[15:0] io_cyclesChannelBusy_292
    //output[15:0] io_cyclesChannelBusy_291
    //output[15:0] io_cyclesChannelBusy_290
    //output[15:0] io_cyclesChannelBusy_289
    //output[15:0] io_cyclesChannelBusy_288
    //output[15:0] io_cyclesChannelBusy_287
    //output[15:0] io_cyclesChannelBusy_286
    //output[15:0] io_cyclesChannelBusy_285
    //output[15:0] io_cyclesChannelBusy_284
    //output[15:0] io_cyclesChannelBusy_283
    //output[15:0] io_cyclesChannelBusy_282
    //output[15:0] io_cyclesChannelBusy_281
    //output[15:0] io_cyclesChannelBusy_280
    //output[15:0] io_cyclesChannelBusy_279
    //output[15:0] io_cyclesChannelBusy_278
    //output[15:0] io_cyclesChannelBusy_277
    //output[15:0] io_cyclesChannelBusy_276
    //output[15:0] io_cyclesChannelBusy_275
    //output[15:0] io_cyclesChannelBusy_274
    //output[15:0] io_cyclesChannelBusy_273
    //output[15:0] io_cyclesChannelBusy_272
    //output[15:0] io_cyclesChannelBusy_271
    //output[15:0] io_cyclesChannelBusy_270
    //output[15:0] io_cyclesChannelBusy_269
    //output[15:0] io_cyclesChannelBusy_268
    //output[15:0] io_cyclesChannelBusy_267
    //output[15:0] io_cyclesChannelBusy_266
    //output[15:0] io_cyclesChannelBusy_265
    //output[15:0] io_cyclesChannelBusy_264
    //output[15:0] io_cyclesChannelBusy_263
    //output[15:0] io_cyclesChannelBusy_262
    //output[15:0] io_cyclesChannelBusy_261
    //output[15:0] io_cyclesChannelBusy_260
    //output[15:0] io_cyclesChannelBusy_259
    //output[15:0] io_cyclesChannelBusy_258
    //output[15:0] io_cyclesChannelBusy_257
    //output[15:0] io_cyclesChannelBusy_256
    //output[15:0] io_cyclesChannelBusy_255
    //output[15:0] io_cyclesChannelBusy_254
    //output[15:0] io_cyclesChannelBusy_253
    //output[15:0] io_cyclesChannelBusy_252
    //output[15:0] io_cyclesChannelBusy_251
    //output[15:0] io_cyclesChannelBusy_250
    //output[15:0] io_cyclesChannelBusy_249
    //output[15:0] io_cyclesChannelBusy_248
    //output[15:0] io_cyclesChannelBusy_247
    //output[15:0] io_cyclesChannelBusy_246
    //output[15:0] io_cyclesChannelBusy_245
    //output[15:0] io_cyclesChannelBusy_244
    //output[15:0] io_cyclesChannelBusy_243
    //output[15:0] io_cyclesChannelBusy_242
    //output[15:0] io_cyclesChannelBusy_241
    //output[15:0] io_cyclesChannelBusy_240
    //output[15:0] io_cyclesChannelBusy_239
    //output[15:0] io_cyclesChannelBusy_238
    //output[15:0] io_cyclesChannelBusy_237
    //output[15:0] io_cyclesChannelBusy_236
    //output[15:0] io_cyclesChannelBusy_235
    //output[15:0] io_cyclesChannelBusy_234
    //output[15:0] io_cyclesChannelBusy_233
    //output[15:0] io_cyclesChannelBusy_232
    //output[15:0] io_cyclesChannelBusy_231
    //output[15:0] io_cyclesChannelBusy_230
    //output[15:0] io_cyclesChannelBusy_229
    //output[15:0] io_cyclesChannelBusy_228
    //output[15:0] io_cyclesChannelBusy_227
    //output[15:0] io_cyclesChannelBusy_226
    //output[15:0] io_cyclesChannelBusy_225
    //output[15:0] io_cyclesChannelBusy_224
    //output[15:0] io_cyclesChannelBusy_223
    //output[15:0] io_cyclesChannelBusy_222
    //output[15:0] io_cyclesChannelBusy_221
    //output[15:0] io_cyclesChannelBusy_220
    //output[15:0] io_cyclesChannelBusy_219
    //output[15:0] io_cyclesChannelBusy_218
    //output[15:0] io_cyclesChannelBusy_217
    //output[15:0] io_cyclesChannelBusy_216
    //output[15:0] io_cyclesChannelBusy_215
    //output[15:0] io_cyclesChannelBusy_214
    //output[15:0] io_cyclesChannelBusy_213
    //output[15:0] io_cyclesChannelBusy_212
    //output[15:0] io_cyclesChannelBusy_211
    //output[15:0] io_cyclesChannelBusy_210
    //output[15:0] io_cyclesChannelBusy_209
    //output[15:0] io_cyclesChannelBusy_208
    //output[15:0] io_cyclesChannelBusy_207
    //output[15:0] io_cyclesChannelBusy_206
    //output[15:0] io_cyclesChannelBusy_205
    //output[15:0] io_cyclesChannelBusy_204
    //output[15:0] io_cyclesChannelBusy_203
    //output[15:0] io_cyclesChannelBusy_202
    //output[15:0] io_cyclesChannelBusy_201
    //output[15:0] io_cyclesChannelBusy_200
    //output[15:0] io_cyclesChannelBusy_199
    //output[15:0] io_cyclesChannelBusy_198
    //output[15:0] io_cyclesChannelBusy_197
    //output[15:0] io_cyclesChannelBusy_196
    //output[15:0] io_cyclesChannelBusy_195
    //output[15:0] io_cyclesChannelBusy_194
    //output[15:0] io_cyclesChannelBusy_193
    //output[15:0] io_cyclesChannelBusy_192
    //output[15:0] io_cyclesChannelBusy_191
    //output[15:0] io_cyclesChannelBusy_190
    //output[15:0] io_cyclesChannelBusy_189
    //output[15:0] io_cyclesChannelBusy_188
    //output[15:0] io_cyclesChannelBusy_187
    //output[15:0] io_cyclesChannelBusy_186
    //output[15:0] io_cyclesChannelBusy_185
    //output[15:0] io_cyclesChannelBusy_184
    //output[15:0] io_cyclesChannelBusy_183
    //output[15:0] io_cyclesChannelBusy_182
    //output[15:0] io_cyclesChannelBusy_181
    //output[15:0] io_cyclesChannelBusy_180
    //output[15:0] io_cyclesChannelBusy_179
    //output[15:0] io_cyclesChannelBusy_178
    //output[15:0] io_cyclesChannelBusy_177
    //output[15:0] io_cyclesChannelBusy_176
    //output[15:0] io_cyclesChannelBusy_175
    //output[15:0] io_cyclesChannelBusy_174
    //output[15:0] io_cyclesChannelBusy_173
    //output[15:0] io_cyclesChannelBusy_172
    //output[15:0] io_cyclesChannelBusy_171
    //output[15:0] io_cyclesChannelBusy_170
    //output[15:0] io_cyclesChannelBusy_169
    //output[15:0] io_cyclesChannelBusy_168
    //output[15:0] io_cyclesChannelBusy_167
    //output[15:0] io_cyclesChannelBusy_166
    //output[15:0] io_cyclesChannelBusy_165
    //output[15:0] io_cyclesChannelBusy_164
    //output[15:0] io_cyclesChannelBusy_163
    //output[15:0] io_cyclesChannelBusy_162
    //output[15:0] io_cyclesChannelBusy_161
    //output[15:0] io_cyclesChannelBusy_160
    //output[15:0] io_cyclesChannelBusy_159
    //output[15:0] io_cyclesChannelBusy_158
    //output[15:0] io_cyclesChannelBusy_157
    //output[15:0] io_cyclesChannelBusy_156
    //output[15:0] io_cyclesChannelBusy_155
    //output[15:0] io_cyclesChannelBusy_154
    //output[15:0] io_cyclesChannelBusy_153
    //output[15:0] io_cyclesChannelBusy_152
    //output[15:0] io_cyclesChannelBusy_151
    //output[15:0] io_cyclesChannelBusy_150
    //output[15:0] io_cyclesChannelBusy_149
    //output[15:0] io_cyclesChannelBusy_148
    //output[15:0] io_cyclesChannelBusy_147
    //output[15:0] io_cyclesChannelBusy_146
    //output[15:0] io_cyclesChannelBusy_145
    //output[15:0] io_cyclesChannelBusy_144
    //output[15:0] io_cyclesChannelBusy_143
    //output[15:0] io_cyclesChannelBusy_142
    //output[15:0] io_cyclesChannelBusy_141
    //output[15:0] io_cyclesChannelBusy_140
    //output[15:0] io_cyclesChannelBusy_139
    //output[15:0] io_cyclesChannelBusy_138
    //output[15:0] io_cyclesChannelBusy_137
    //output[15:0] io_cyclesChannelBusy_136
    //output[15:0] io_cyclesChannelBusy_135
    //output[15:0] io_cyclesChannelBusy_134
    //output[15:0] io_cyclesChannelBusy_133
    //output[15:0] io_cyclesChannelBusy_132
    //output[15:0] io_cyclesChannelBusy_131
    //output[15:0] io_cyclesChannelBusy_130
    //output[15:0] io_cyclesChannelBusy_129
    //output[15:0] io_cyclesChannelBusy_128
    //output[15:0] io_cyclesChannelBusy_127
    //output[15:0] io_cyclesChannelBusy_126
    //output[15:0] io_cyclesChannelBusy_125
    //output[15:0] io_cyclesChannelBusy_124
    //output[15:0] io_cyclesChannelBusy_123
    //output[15:0] io_cyclesChannelBusy_122
    //output[15:0] io_cyclesChannelBusy_121
    //output[15:0] io_cyclesChannelBusy_120
    //output[15:0] io_cyclesChannelBusy_119
    //output[15:0] io_cyclesChannelBusy_118
    //output[15:0] io_cyclesChannelBusy_117
    //output[15:0] io_cyclesChannelBusy_116
    //output[15:0] io_cyclesChannelBusy_115
    //output[15:0] io_cyclesChannelBusy_114
    //output[15:0] io_cyclesChannelBusy_113
    //output[15:0] io_cyclesChannelBusy_112
    //output[15:0] io_cyclesChannelBusy_111
    //output[15:0] io_cyclesChannelBusy_110
    //output[15:0] io_cyclesChannelBusy_109
    //output[15:0] io_cyclesChannelBusy_108
    //output[15:0] io_cyclesChannelBusy_107
    //output[15:0] io_cyclesChannelBusy_106
    //output[15:0] io_cyclesChannelBusy_105
    //output[15:0] io_cyclesChannelBusy_104
    //output[15:0] io_cyclesChannelBusy_103
    //output[15:0] io_cyclesChannelBusy_102
    //output[15:0] io_cyclesChannelBusy_101
    //output[15:0] io_cyclesChannelBusy_100
    //output[15:0] io_cyclesChannelBusy_99
    //output[15:0] io_cyclesChannelBusy_98
    //output[15:0] io_cyclesChannelBusy_97
    //output[15:0] io_cyclesChannelBusy_96
    //output[15:0] io_cyclesChannelBusy_95
    //output[15:0] io_cyclesChannelBusy_94
    //output[15:0] io_cyclesChannelBusy_93
    //output[15:0] io_cyclesChannelBusy_92
    //output[15:0] io_cyclesChannelBusy_91
    //output[15:0] io_cyclesChannelBusy_90
    //output[15:0] io_cyclesChannelBusy_89
    //output[15:0] io_cyclesChannelBusy_88
    //output[15:0] io_cyclesChannelBusy_87
    //output[15:0] io_cyclesChannelBusy_86
    //output[15:0] io_cyclesChannelBusy_85
    //output[15:0] io_cyclesChannelBusy_84
    //output[15:0] io_cyclesChannelBusy_83
    //output[15:0] io_cyclesChannelBusy_82
    //output[15:0] io_cyclesChannelBusy_81
    //output[15:0] io_cyclesChannelBusy_80
    //output[15:0] io_cyclesChannelBusy_79
    //output[15:0] io_cyclesChannelBusy_78
    //output[15:0] io_cyclesChannelBusy_77
    //output[15:0] io_cyclesChannelBusy_76
    //output[15:0] io_cyclesChannelBusy_75
    //output[15:0] io_cyclesChannelBusy_74
    //output[15:0] io_cyclesChannelBusy_73
    //output[15:0] io_cyclesChannelBusy_72
    //output[15:0] io_cyclesChannelBusy_71
    //output[15:0] io_cyclesChannelBusy_70
    //output[15:0] io_cyclesChannelBusy_69
    //output[15:0] io_cyclesChannelBusy_68
    //output[15:0] io_cyclesChannelBusy_67
    //output[15:0] io_cyclesChannelBusy_66
    //output[15:0] io_cyclesChannelBusy_65
    //output[15:0] io_cyclesChannelBusy_64
    //output[15:0] io_cyclesChannelBusy_63
    //output[15:0] io_cyclesChannelBusy_62
    //output[15:0] io_cyclesChannelBusy_61
    //output[15:0] io_cyclesChannelBusy_60
    //output[15:0] io_cyclesChannelBusy_59
    //output[15:0] io_cyclesChannelBusy_58
    //output[15:0] io_cyclesChannelBusy_57
    //output[15:0] io_cyclesChannelBusy_56
    //output[15:0] io_cyclesChannelBusy_55
    //output[15:0] io_cyclesChannelBusy_54
    //output[15:0] io_cyclesChannelBusy_53
    //output[15:0] io_cyclesChannelBusy_52
    //output[15:0] io_cyclesChannelBusy_51
    //output[15:0] io_cyclesChannelBusy_50
    //output[15:0] io_cyclesChannelBusy_49
    //output[15:0] io_cyclesChannelBusy_48
    //output[15:0] io_cyclesChannelBusy_47
    //output[15:0] io_cyclesChannelBusy_46
    //output[15:0] io_cyclesChannelBusy_45
    //output[15:0] io_cyclesChannelBusy_44
    //output[15:0] io_cyclesChannelBusy_43
    //output[15:0] io_cyclesChannelBusy_42
    //output[15:0] io_cyclesChannelBusy_41
    //output[15:0] io_cyclesChannelBusy_40
    //output[15:0] io_cyclesChannelBusy_39
    //output[15:0] io_cyclesChannelBusy_38
    //output[15:0] io_cyclesChannelBusy_37
    //output[15:0] io_cyclesChannelBusy_36
    //output[15:0] io_cyclesChannelBusy_35
    //output[15:0] io_cyclesChannelBusy_34
    //output[15:0] io_cyclesChannelBusy_33
    //output[15:0] io_cyclesChannelBusy_32
    //output[15:0] io_cyclesChannelBusy_31
    //output[15:0] io_cyclesChannelBusy_30
    //output[15:0] io_cyclesChannelBusy_29
    //output[15:0] io_cyclesChannelBusy_28
    //output[15:0] io_cyclesChannelBusy_27
    //output[15:0] io_cyclesChannelBusy_26
    //output[15:0] io_cyclesChannelBusy_25
    //output[15:0] io_cyclesChannelBusy_24
    //output[15:0] io_cyclesChannelBusy_23
    //output[15:0] io_cyclesChannelBusy_22
    //output[15:0] io_cyclesChannelBusy_21
    //output[15:0] io_cyclesChannelBusy_20
    //output[15:0] io_cyclesChannelBusy_19
    //output[15:0] io_cyclesChannelBusy_18
    //output[15:0] io_cyclesChannelBusy_17
    //output[15:0] io_cyclesChannelBusy_16
    //output[15:0] io_cyclesChannelBusy_15
    output[15:0] io_cyclesChannelBusy_14,
    output[15:0] io_cyclesChannelBusy_13,
    output[15:0] io_cyclesChannelBusy_12,
    output[15:0] io_cyclesChannelBusy_11,
    output[15:0] io_cyclesChannelBusy_10,
    output[15:0] io_cyclesChannelBusy_9,
    output[15:0] io_cyclesChannelBusy_8,
    output[15:0] io_cyclesChannelBusy_7,
    output[15:0] io_cyclesChannelBusy_6,
    output[15:0] io_cyclesChannelBusy_5,
    output[15:0] io_cyclesChannelBusy_4,
    output[15:0] io_cyclesChannelBusy_3,
    output[15:0] io_cyclesChannelBusy_2,
    output[15:0] io_cyclesChannelBusy_1,
    output[15:0] io_cyclesChannelBusy_0,
    input  io_bypass_2,
    input  io_bypass_1,
    input  io_bypass_0
);

  wire[15:0] BusProbe_io_cyclesChannelBusy_1;
  wire[15:0] BusProbe_io_cyclesRouterBusy;
  wire CreditBuffer_io_in_1_credit_1_grant;
  wire CreditBuffer_io_in_1_credit_0_grant;
  wire[54:0] CreditBuffer_io_out_1_flit_x;
  wire CreditBuffer_io_out_1_flitValid;
  wire[15:0] BusProbe_1_io_cyclesChannelBusy_2;
  wire[15:0] BusProbe_1_io_cyclesChannelBusy_1;
  wire[15:0] BusProbe_1_io_cyclesRouterBusy;
  wire CreditBuffer_1_io_in_2_credit_1_grant;
  wire CreditBuffer_1_io_in_2_credit_0_grant;
  wire CreditBuffer_1_io_in_1_credit_1_grant;
  wire CreditBuffer_1_io_in_1_credit_0_grant;
  wire[54:0] CreditBuffer_1_io_out_2_flit_x;
  wire CreditBuffer_1_io_out_2_flitValid;
  wire[54:0] CreditBuffer_1_io_out_1_flit_x;
  wire CreditBuffer_1_io_out_1_flitValid;
  wire[15:0] BusProbe_2_io_cyclesChannelBusy_2;
  wire[15:0] BusProbe_2_io_cyclesRouterBusy;
  wire CreditBuffer_2_io_in_2_credit_1_grant;
  wire CreditBuffer_2_io_in_2_credit_0_grant;
  wire[54:0] CreditBuffer_2_io_out_2_flit_x;
  wire CreditBuffer_2_io_out_2_flitValid;
  wire[54:0] OpenSoC_VCConstantEndpoint_io_outChannels_1_flit_x;
  wire OpenSoC_VCConstantEndpoint_io_outChannels_1_flitValid;
  wire[54:0] OpenSoC_VCConstantEndpoint_1_io_outChannels_3_flit_x;
  wire OpenSoC_VCConstantEndpoint_1_io_outChannels_3_flitValid;
  wire[54:0] OpenSoC_VCConstantEndpoint_2_io_outChannels_4_flit_x;
  wire OpenSoC_VCConstantEndpoint_2_io_outChannels_4_flitValid;
  wire[54:0] OpenSoC_VCConstantEndpoint_3_io_outChannels_3_flit_x;
  wire OpenSoC_VCConstantEndpoint_3_io_outChannels_3_flitValid;
  wire[54:0] OpenSoC_VCConstantEndpoint_4_io_outChannels_4_flit_x;
  wire OpenSoC_VCConstantEndpoint_4_io_outChannels_4_flitValid;
  wire[54:0] OpenSoC_VCConstantEndpoint_5_io_outChannels_2_flit_x;
  wire OpenSoC_VCConstantEndpoint_5_io_outChannels_2_flitValid;
  wire[54:0] OpenSoC_VCConstantEndpoint_6_io_outChannels_3_flit_x;
  wire OpenSoC_VCConstantEndpoint_6_io_outChannels_3_flitValid;
  wire[54:0] OpenSoC_VCConstantEndpoint_7_io_outChannels_4_flit_x;
  wire OpenSoC_VCConstantEndpoint_7_io_outChannels_4_flitValid;
  wire VCRouterWrapper_io_inChannels_4_credit_1_grant;
  wire VCRouterWrapper_io_inChannels_4_credit_0_grant;
  wire VCRouterWrapper_io_inChannels_3_credit_1_grant;
  wire VCRouterWrapper_io_inChannels_3_credit_0_grant;
  wire VCRouterWrapper_io_inChannels_2_credit_1_grant;
  wire VCRouterWrapper_io_inChannels_2_credit_0_grant;
  wire VCRouterWrapper_io_inChannels_1_credit_1_grant;
  wire VCRouterWrapper_io_inChannels_1_credit_0_grant;
  wire VCRouterWrapper_io_inChannels_0_credit_1_grant;
  wire VCRouterWrapper_io_inChannels_0_credit_0_grant;
  wire[54:0] VCRouterWrapper_io_outChannels_4_flit_x;
  wire VCRouterWrapper_io_outChannels_4_flitValid;
  wire[54:0] VCRouterWrapper_io_outChannels_3_flit_x;
  wire VCRouterWrapper_io_outChannels_3_flitValid;
  wire[54:0] VCRouterWrapper_io_outChannels_1_flit_x;
  wire VCRouterWrapper_io_outChannels_1_flitValid;
  wire[54:0] VCRouterWrapper_io_outChannels_0_flit_x;
  wire VCRouterWrapper_io_outChannels_0_flitValid;
  wire VCRouterWrapper_1_io_inChannels_4_credit_1_grant;
  wire VCRouterWrapper_1_io_inChannels_4_credit_0_grant;
  wire VCRouterWrapper_1_io_inChannels_3_credit_1_grant;
  wire VCRouterWrapper_1_io_inChannels_3_credit_0_grant;
  wire VCRouterWrapper_1_io_inChannels_2_credit_1_grant;
  wire VCRouterWrapper_1_io_inChannels_2_credit_0_grant;
  wire VCRouterWrapper_1_io_inChannels_1_credit_1_grant;
  wire VCRouterWrapper_1_io_inChannels_1_credit_0_grant;
  wire VCRouterWrapper_1_io_inChannels_0_credit_1_grant;
  wire VCRouterWrapper_1_io_inChannels_0_credit_0_grant;
  wire[54:0] VCRouterWrapper_1_io_outChannels_4_flit_x;
  wire VCRouterWrapper_1_io_outChannels_4_flitValid;
  wire[54:0] VCRouterWrapper_1_io_outChannels_3_flit_x;
  wire VCRouterWrapper_1_io_outChannels_3_flitValid;
  wire[54:0] VCRouterWrapper_1_io_outChannels_2_flit_x;
  wire VCRouterWrapper_1_io_outChannels_2_flitValid;
  wire[54:0] VCRouterWrapper_1_io_outChannels_1_flit_x;
  wire VCRouterWrapper_1_io_outChannels_1_flitValid;
  wire[54:0] VCRouterWrapper_1_io_outChannels_0_flit_x;
  wire VCRouterWrapper_1_io_outChannels_0_flitValid;
  wire VCRouterWrapper_2_io_inChannels_4_credit_1_grant;
  wire VCRouterWrapper_2_io_inChannels_4_credit_0_grant;
  wire VCRouterWrapper_2_io_inChannels_3_credit_1_grant;
  wire VCRouterWrapper_2_io_inChannels_3_credit_0_grant;
  wire VCRouterWrapper_2_io_inChannels_2_credit_1_grant;
  wire VCRouterWrapper_2_io_inChannels_2_credit_0_grant;
  wire VCRouterWrapper_2_io_inChannels_1_credit_1_grant;
  wire VCRouterWrapper_2_io_inChannels_1_credit_0_grant;
  wire VCRouterWrapper_2_io_inChannels_0_credit_1_grant;
  wire VCRouterWrapper_2_io_inChannels_0_credit_0_grant;
  wire[54:0] VCRouterWrapper_2_io_outChannels_4_flit_x;
  wire VCRouterWrapper_2_io_outChannels_4_flitValid;
  wire[54:0] VCRouterWrapper_2_io_outChannels_3_flit_x;
  wire VCRouterWrapper_2_io_outChannels_3_flitValid;
  wire[54:0] VCRouterWrapper_2_io_outChannels_2_flit_x;
  wire VCRouterWrapper_2_io_outChannels_2_flitValid;
  wire[54:0] VCRouterWrapper_2_io_outChannels_0_flit_x;
  wire VCRouterWrapper_2_io_outChannels_0_flitValid;


`ifndef SYNTHESIS
// synthesis translate_off
  assign io_cyclesChannelBusy_0 = {1{1'b0}};
  assign io_cyclesChannelBusy_2 = {1{1'b0}};
  assign io_cyclesChannelBusy_3 = {1{1'b0}};
  assign io_cyclesChannelBusy_4 = {1{1'b0}};
  assign io_cyclesChannelBusy_5 = {1{1'b0}};
  assign io_cyclesChannelBusy_8 = {1{1'b0}};
  assign io_cyclesChannelBusy_9 = {1{1'b0}};
  assign io_cyclesChannelBusy_10 = {1{1'b0}};
  assign io_cyclesChannelBusy_11 = {1{1'b0}};
  assign io_cyclesChannelBusy_13 = {1{1'b0}};
  assign io_cyclesChannelBusy_14 = {1{1'b0}};
//  assign io_cyclesChannelBusy_15 = {1{1'b0}};
//  assign io_cyclesChannelBusy_16 = {1{1'b0}};
//  assign io_cyclesChannelBusy_17 = {1{1'b0}};
//  assign io_cyclesChannelBusy_18 = {1{1'b0}};
//  assign io_cyclesChannelBusy_19 = {1{1'b0}};
//  assign io_cyclesChannelBusy_20 = {1{1'b0}};
//  assign io_cyclesChannelBusy_21 = {1{1'b0}};
//  assign io_cyclesChannelBusy_22 = {1{1'b0}};
//  assign io_cyclesChannelBusy_23 = {1{1'b0}};
//  assign io_cyclesChannelBusy_24 = {1{1'b0}};
//  assign io_cyclesChannelBusy_25 = {1{1'b0}};
//  assign io_cyclesChannelBusy_26 = {1{1'b0}};
//  assign io_cyclesChannelBusy_27 = {1{1'b0}};
//  assign io_cyclesChannelBusy_28 = {1{1'b0}};
//  assign io_cyclesChannelBusy_29 = {1{1'b0}};
//  assign io_cyclesChannelBusy_30 = {1{1'b0}};
//  assign io_cyclesChannelBusy_31 = {1{1'b0}};
//  assign io_cyclesChannelBusy_32 = {1{1'b0}};
//  assign io_cyclesChannelBusy_33 = {1{1'b0}};
//  assign io_cyclesChannelBusy_34 = {1{1'b0}};
//  assign io_cyclesChannelBusy_35 = {1{1'b0}};
//  assign io_cyclesChannelBusy_36 = {1{1'b0}};
//  assign io_cyclesChannelBusy_37 = {1{1'b0}};
//  assign io_cyclesChannelBusy_38 = {1{1'b0}};
//  assign io_cyclesChannelBusy_39 = {1{1'b0}};
//  assign io_cyclesChannelBusy_40 = {1{1'b0}};
//  assign io_cyclesChannelBusy_41 = {1{1'b0}};
//  assign io_cyclesChannelBusy_42 = {1{1'b0}};
//  assign io_cyclesChannelBusy_43 = {1{1'b0}};
//  assign io_cyclesChannelBusy_44 = {1{1'b0}};
//  assign io_cyclesChannelBusy_45 = {1{1'b0}};
//  assign io_cyclesChannelBusy_46 = {1{1'b0}};
//  assign io_cyclesChannelBusy_47 = {1{1'b0}};
//  assign io_cyclesChannelBusy_48 = {1{1'b0}};
//  assign io_cyclesChannelBusy_49 = {1{1'b0}};
//  assign io_cyclesChannelBusy_50 = {1{1'b0}};
//  assign io_cyclesChannelBusy_51 = {1{1'b0}};
//  assign io_cyclesChannelBusy_52 = {1{1'b0}};
//  assign io_cyclesChannelBusy_53 = {1{1'b0}};
//  assign io_cyclesChannelBusy_54 = {1{1'b0}};
//  assign io_cyclesChannelBusy_55 = {1{1'b0}};
//  assign io_cyclesChannelBusy_56 = {1{1'b0}};
//  assign io_cyclesChannelBusy_57 = {1{1'b0}};
//  assign io_cyclesChannelBusy_58 = {1{1'b0}};
//  assign io_cyclesChannelBusy_59 = {1{1'b0}};
//  assign io_cyclesChannelBusy_60 = {1{1'b0}};
//  assign io_cyclesChannelBusy_61 = {1{1'b0}};
//  assign io_cyclesChannelBusy_62 = {1{1'b0}};
//  assign io_cyclesChannelBusy_63 = {1{1'b0}};
//  assign io_cyclesChannelBusy_64 = {1{1'b0}};
//  assign io_cyclesChannelBusy_65 = {1{1'b0}};
//  assign io_cyclesChannelBusy_66 = {1{1'b0}};
//  assign io_cyclesChannelBusy_67 = {1{1'b0}};
//  assign io_cyclesChannelBusy_68 = {1{1'b0}};
//  assign io_cyclesChannelBusy_69 = {1{1'b0}};
//  assign io_cyclesChannelBusy_70 = {1{1'b0}};
//  assign io_cyclesChannelBusy_71 = {1{1'b0}};
//  assign io_cyclesChannelBusy_72 = {1{1'b0}};
//  assign io_cyclesChannelBusy_73 = {1{1'b0}};
//  assign io_cyclesChannelBusy_74 = {1{1'b0}};
//  assign io_cyclesChannelBusy_75 = {1{1'b0}};
//  assign io_cyclesChannelBusy_76 = {1{1'b0}};
//  assign io_cyclesChannelBusy_77 = {1{1'b0}};
//  assign io_cyclesChannelBusy_78 = {1{1'b0}};
//  assign io_cyclesChannelBusy_79 = {1{1'b0}};
//  assign io_cyclesChannelBusy_80 = {1{1'b0}};
//  assign io_cyclesChannelBusy_81 = {1{1'b0}};
//  assign io_cyclesChannelBusy_82 = {1{1'b0}};
//  assign io_cyclesChannelBusy_83 = {1{1'b0}};
//  assign io_cyclesChannelBusy_84 = {1{1'b0}};
//  assign io_cyclesChannelBusy_85 = {1{1'b0}};
//  assign io_cyclesChannelBusy_86 = {1{1'b0}};
//  assign io_cyclesChannelBusy_87 = {1{1'b0}};
//  assign io_cyclesChannelBusy_88 = {1{1'b0}};
//  assign io_cyclesChannelBusy_89 = {1{1'b0}};
//  assign io_cyclesChannelBusy_90 = {1{1'b0}};
//  assign io_cyclesChannelBusy_91 = {1{1'b0}};
//  assign io_cyclesChannelBusy_92 = {1{1'b0}};
//  assign io_cyclesChannelBusy_93 = {1{1'b0}};
//  assign io_cyclesChannelBusy_94 = {1{1'b0}};
//  assign io_cyclesChannelBusy_95 = {1{1'b0}};
//  assign io_cyclesChannelBusy_96 = {1{1'b0}};
//  assign io_cyclesChannelBusy_97 = {1{1'b0}};
//  assign io_cyclesChannelBusy_98 = {1{1'b0}};
//  assign io_cyclesChannelBusy_99 = {1{1'b0}};
//  assign io_cyclesChannelBusy_100 = {1{1'b0}};
//  assign io_cyclesChannelBusy_101 = {1{1'b0}};
//  assign io_cyclesChannelBusy_102 = {1{1'b0}};
//  assign io_cyclesChannelBusy_103 = {1{1'b0}};
//  assign io_cyclesChannelBusy_104 = {1{1'b0}};
//  assign io_cyclesChannelBusy_105 = {1{1'b0}};
//  assign io_cyclesChannelBusy_106 = {1{1'b0}};
//  assign io_cyclesChannelBusy_107 = {1{1'b0}};
//  assign io_cyclesChannelBusy_108 = {1{1'b0}};
//  assign io_cyclesChannelBusy_109 = {1{1'b0}};
//  assign io_cyclesChannelBusy_110 = {1{1'b0}};
//  assign io_cyclesChannelBusy_111 = {1{1'b0}};
//  assign io_cyclesChannelBusy_112 = {1{1'b0}};
//  assign io_cyclesChannelBusy_113 = {1{1'b0}};
//  assign io_cyclesChannelBusy_114 = {1{1'b0}};
//  assign io_cyclesChannelBusy_115 = {1{1'b0}};
//  assign io_cyclesChannelBusy_116 = {1{1'b0}};
//  assign io_cyclesChannelBusy_117 = {1{1'b0}};
//  assign io_cyclesChannelBusy_118 = {1{1'b0}};
//  assign io_cyclesChannelBusy_119 = {1{1'b0}};
//  assign io_cyclesChannelBusy_120 = {1{1'b0}};
//  assign io_cyclesChannelBusy_121 = {1{1'b0}};
//  assign io_cyclesChannelBusy_122 = {1{1'b0}};
//  assign io_cyclesChannelBusy_123 = {1{1'b0}};
//  assign io_cyclesChannelBusy_124 = {1{1'b0}};
//  assign io_cyclesChannelBusy_125 = {1{1'b0}};
//  assign io_cyclesChannelBusy_126 = {1{1'b0}};
//  assign io_cyclesChannelBusy_127 = {1{1'b0}};
//  assign io_cyclesChannelBusy_128 = {1{1'b0}};
//  assign io_cyclesChannelBusy_129 = {1{1'b0}};
//  assign io_cyclesChannelBusy_130 = {1{1'b0}};
//  assign io_cyclesChannelBusy_131 = {1{1'b0}};
//  assign io_cyclesChannelBusy_132 = {1{1'b0}};
//  assign io_cyclesChannelBusy_133 = {1{1'b0}};
//  assign io_cyclesChannelBusy_134 = {1{1'b0}};
//  assign io_cyclesChannelBusy_135 = {1{1'b0}};
//  assign io_cyclesChannelBusy_136 = {1{1'b0}};
//  assign io_cyclesChannelBusy_137 = {1{1'b0}};
//  assign io_cyclesChannelBusy_138 = {1{1'b0}};
//  assign io_cyclesChannelBusy_139 = {1{1'b0}};
//  assign io_cyclesChannelBusy_140 = {1{1'b0}};
//  assign io_cyclesChannelBusy_141 = {1{1'b0}};
//  assign io_cyclesChannelBusy_142 = {1{1'b0}};
//  assign io_cyclesChannelBusy_143 = {1{1'b0}};
//  assign io_cyclesChannelBusy_144 = {1{1'b0}};
//  assign io_cyclesChannelBusy_145 = {1{1'b0}};
//  assign io_cyclesChannelBusy_146 = {1{1'b0}};
//  assign io_cyclesChannelBusy_147 = {1{1'b0}};
//  assign io_cyclesChannelBusy_148 = {1{1'b0}};
//  assign io_cyclesChannelBusy_149 = {1{1'b0}};
//  assign io_cyclesChannelBusy_150 = {1{1'b0}};
//  assign io_cyclesChannelBusy_151 = {1{1'b0}};
//  assign io_cyclesChannelBusy_152 = {1{1'b0}};
//  assign io_cyclesChannelBusy_153 = {1{1'b0}};
//  assign io_cyclesChannelBusy_154 = {1{1'b0}};
//  assign io_cyclesChannelBusy_155 = {1{1'b0}};
//  assign io_cyclesChannelBusy_156 = {1{1'b0}};
//  assign io_cyclesChannelBusy_157 = {1{1'b0}};
//  assign io_cyclesChannelBusy_158 = {1{1'b0}};
//  assign io_cyclesChannelBusy_159 = {1{1'b0}};
//  assign io_cyclesChannelBusy_160 = {1{1'b0}};
//  assign io_cyclesChannelBusy_161 = {1{1'b0}};
//  assign io_cyclesChannelBusy_162 = {1{1'b0}};
//  assign io_cyclesChannelBusy_163 = {1{1'b0}};
//  assign io_cyclesChannelBusy_164 = {1{1'b0}};
//  assign io_cyclesChannelBusy_165 = {1{1'b0}};
//  assign io_cyclesChannelBusy_166 = {1{1'b0}};
//  assign io_cyclesChannelBusy_167 = {1{1'b0}};
//  assign io_cyclesChannelBusy_168 = {1{1'b0}};
//  assign io_cyclesChannelBusy_169 = {1{1'b0}};
//  assign io_cyclesChannelBusy_170 = {1{1'b0}};
//  assign io_cyclesChannelBusy_171 = {1{1'b0}};
//  assign io_cyclesChannelBusy_172 = {1{1'b0}};
//  assign io_cyclesChannelBusy_173 = {1{1'b0}};
//  assign io_cyclesChannelBusy_174 = {1{1'b0}};
//  assign io_cyclesChannelBusy_175 = {1{1'b0}};
//  assign io_cyclesChannelBusy_176 = {1{1'b0}};
//  assign io_cyclesChannelBusy_177 = {1{1'b0}};
//  assign io_cyclesChannelBusy_178 = {1{1'b0}};
//  assign io_cyclesChannelBusy_179 = {1{1'b0}};
//  assign io_cyclesChannelBusy_180 = {1{1'b0}};
//  assign io_cyclesChannelBusy_181 = {1{1'b0}};
//  assign io_cyclesChannelBusy_182 = {1{1'b0}};
//  assign io_cyclesChannelBusy_183 = {1{1'b0}};
//  assign io_cyclesChannelBusy_184 = {1{1'b0}};
//  assign io_cyclesChannelBusy_185 = {1{1'b0}};
//  assign io_cyclesChannelBusy_186 = {1{1'b0}};
//  assign io_cyclesChannelBusy_187 = {1{1'b0}};
//  assign io_cyclesChannelBusy_188 = {1{1'b0}};
//  assign io_cyclesChannelBusy_189 = {1{1'b0}};
//  assign io_cyclesChannelBusy_190 = {1{1'b0}};
//  assign io_cyclesChannelBusy_191 = {1{1'b0}};
//  assign io_cyclesChannelBusy_192 = {1{1'b0}};
//  assign io_cyclesChannelBusy_193 = {1{1'b0}};
//  assign io_cyclesChannelBusy_194 = {1{1'b0}};
//  assign io_cyclesChannelBusy_195 = {1{1'b0}};
//  assign io_cyclesChannelBusy_196 = {1{1'b0}};
//  assign io_cyclesChannelBusy_197 = {1{1'b0}};
//  assign io_cyclesChannelBusy_198 = {1{1'b0}};
//  assign io_cyclesChannelBusy_199 = {1{1'b0}};
//  assign io_cyclesChannelBusy_200 = {1{1'b0}};
//  assign io_cyclesChannelBusy_201 = {1{1'b0}};
//  assign io_cyclesChannelBusy_202 = {1{1'b0}};
//  assign io_cyclesChannelBusy_203 = {1{1'b0}};
//  assign io_cyclesChannelBusy_204 = {1{1'b0}};
//  assign io_cyclesChannelBusy_205 = {1{1'b0}};
//  assign io_cyclesChannelBusy_206 = {1{1'b0}};
//  assign io_cyclesChannelBusy_207 = {1{1'b0}};
//  assign io_cyclesChannelBusy_208 = {1{1'b0}};
//  assign io_cyclesChannelBusy_209 = {1{1'b0}};
//  assign io_cyclesChannelBusy_210 = {1{1'b0}};
//  assign io_cyclesChannelBusy_211 = {1{1'b0}};
//  assign io_cyclesChannelBusy_212 = {1{1'b0}};
//  assign io_cyclesChannelBusy_213 = {1{1'b0}};
//  assign io_cyclesChannelBusy_214 = {1{1'b0}};
//  assign io_cyclesChannelBusy_215 = {1{1'b0}};
//  assign io_cyclesChannelBusy_216 = {1{1'b0}};
//  assign io_cyclesChannelBusy_217 = {1{1'b0}};
//  assign io_cyclesChannelBusy_218 = {1{1'b0}};
//  assign io_cyclesChannelBusy_219 = {1{1'b0}};
//  assign io_cyclesChannelBusy_220 = {1{1'b0}};
//  assign io_cyclesChannelBusy_221 = {1{1'b0}};
//  assign io_cyclesChannelBusy_222 = {1{1'b0}};
//  assign io_cyclesChannelBusy_223 = {1{1'b0}};
//  assign io_cyclesChannelBusy_224 = {1{1'b0}};
//  assign io_cyclesChannelBusy_225 = {1{1'b0}};
//  assign io_cyclesChannelBusy_226 = {1{1'b0}};
//  assign io_cyclesChannelBusy_227 = {1{1'b0}};
//  assign io_cyclesChannelBusy_228 = {1{1'b0}};
//  assign io_cyclesChannelBusy_229 = {1{1'b0}};
//  assign io_cyclesChannelBusy_230 = {1{1'b0}};
//  assign io_cyclesChannelBusy_231 = {1{1'b0}};
//  assign io_cyclesChannelBusy_232 = {1{1'b0}};
//  assign io_cyclesChannelBusy_233 = {1{1'b0}};
//  assign io_cyclesChannelBusy_234 = {1{1'b0}};
//  assign io_cyclesChannelBusy_235 = {1{1'b0}};
//  assign io_cyclesChannelBusy_236 = {1{1'b0}};
//  assign io_cyclesChannelBusy_237 = {1{1'b0}};
//  assign io_cyclesChannelBusy_238 = {1{1'b0}};
//  assign io_cyclesChannelBusy_239 = {1{1'b0}};
//  assign io_cyclesChannelBusy_240 = {1{1'b0}};
//  assign io_cyclesChannelBusy_241 = {1{1'b0}};
//  assign io_cyclesChannelBusy_242 = {1{1'b0}};
//  assign io_cyclesChannelBusy_243 = {1{1'b0}};
//  assign io_cyclesChannelBusy_244 = {1{1'b0}};
//  assign io_cyclesChannelBusy_245 = {1{1'b0}};
//  assign io_cyclesChannelBusy_246 = {1{1'b0}};
//  assign io_cyclesChannelBusy_247 = {1{1'b0}};
//  assign io_cyclesChannelBusy_248 = {1{1'b0}};
//  assign io_cyclesChannelBusy_249 = {1{1'b0}};
//  assign io_cyclesChannelBusy_250 = {1{1'b0}};
//  assign io_cyclesChannelBusy_251 = {1{1'b0}};
//  assign io_cyclesChannelBusy_252 = {1{1'b0}};
//  assign io_cyclesChannelBusy_253 = {1{1'b0}};
//  assign io_cyclesChannelBusy_254 = {1{1'b0}};
//  assign io_cyclesChannelBusy_255 = {1{1'b0}};
//  assign io_cyclesChannelBusy_256 = {1{1'b0}};
//  assign io_cyclesChannelBusy_257 = {1{1'b0}};
//  assign io_cyclesChannelBusy_258 = {1{1'b0}};
//  assign io_cyclesChannelBusy_259 = {1{1'b0}};
//  assign io_cyclesChannelBusy_260 = {1{1'b0}};
//  assign io_cyclesChannelBusy_261 = {1{1'b0}};
//  assign io_cyclesChannelBusy_262 = {1{1'b0}};
//  assign io_cyclesChannelBusy_263 = {1{1'b0}};
//  assign io_cyclesChannelBusy_264 = {1{1'b0}};
//  assign io_cyclesChannelBusy_265 = {1{1'b0}};
//  assign io_cyclesChannelBusy_266 = {1{1'b0}};
//  assign io_cyclesChannelBusy_267 = {1{1'b0}};
//  assign io_cyclesChannelBusy_268 = {1{1'b0}};
//  assign io_cyclesChannelBusy_269 = {1{1'b0}};
//  assign io_cyclesChannelBusy_270 = {1{1'b0}};
//  assign io_cyclesChannelBusy_271 = {1{1'b0}};
//  assign io_cyclesChannelBusy_272 = {1{1'b0}};
//  assign io_cyclesChannelBusy_273 = {1{1'b0}};
//  assign io_cyclesChannelBusy_274 = {1{1'b0}};
//  assign io_cyclesChannelBusy_275 = {1{1'b0}};
//  assign io_cyclesChannelBusy_276 = {1{1'b0}};
//  assign io_cyclesChannelBusy_277 = {1{1'b0}};
//  assign io_cyclesChannelBusy_278 = {1{1'b0}};
//  assign io_cyclesChannelBusy_279 = {1{1'b0}};
//  assign io_cyclesChannelBusy_280 = {1{1'b0}};
//  assign io_cyclesChannelBusy_281 = {1{1'b0}};
//  assign io_cyclesChannelBusy_282 = {1{1'b0}};
//  assign io_cyclesChannelBusy_283 = {1{1'b0}};
//  assign io_cyclesChannelBusy_284 = {1{1'b0}};
//  assign io_cyclesChannelBusy_285 = {1{1'b0}};
//  assign io_cyclesChannelBusy_286 = {1{1'b0}};
//  assign io_cyclesChannelBusy_287 = {1{1'b0}};
//  assign io_cyclesChannelBusy_288 = {1{1'b0}};
//  assign io_cyclesChannelBusy_289 = {1{1'b0}};
//  assign io_cyclesChannelBusy_290 = {1{1'b0}};
//  assign io_cyclesChannelBusy_291 = {1{1'b0}};
//  assign io_cyclesChannelBusy_292 = {1{1'b0}};
//  assign io_cyclesChannelBusy_293 = {1{1'b0}};
//  assign io_cyclesChannelBusy_294 = {1{1'b0}};
//  assign io_cyclesChannelBusy_295 = {1{1'b0}};
//  assign io_cyclesChannelBusy_296 = {1{1'b0}};
//  assign io_cyclesChannelBusy_297 = {1{1'b0}};
//  assign io_cyclesChannelBusy_298 = {1{1'b0}};
//  assign io_cyclesChannelBusy_299 = {1{1'b0}};
//  assign io_cyclesChannelBusy_300 = {1{1'b0}};
//  assign io_cyclesChannelBusy_301 = {1{1'b0}};
//  assign io_cyclesChannelBusy_302 = {1{1'b0}};
//  assign io_cyclesChannelBusy_303 = {1{1'b0}};
//  assign io_cyclesChannelBusy_304 = {1{1'b0}};
//  assign io_cyclesChannelBusy_305 = {1{1'b0}};
//  assign io_cyclesChannelBusy_306 = {1{1'b0}};
//  assign io_cyclesChannelBusy_307 = {1{1'b0}};
//  assign io_cyclesChannelBusy_308 = {1{1'b0}};
//  assign io_cyclesChannelBusy_309 = {1{1'b0}};
//  assign io_cyclesChannelBusy_310 = {1{1'b0}};
//  assign io_cyclesChannelBusy_311 = {1{1'b0}};
//  assign io_cyclesChannelBusy_312 = {1{1'b0}};
//  assign io_cyclesChannelBusy_313 = {1{1'b0}};
//  assign io_cyclesChannelBusy_314 = {1{1'b0}};
//  assign io_cyclesChannelBusy_315 = {1{1'b0}};
//  assign io_cyclesChannelBusy_316 = {1{1'b0}};
//  assign io_cyclesChannelBusy_317 = {1{1'b0}};
//  assign io_cyclesChannelBusy_318 = {1{1'b0}};
//  assign io_cyclesChannelBusy_319 = {1{1'b0}};
//  assign io_cyclesChannelBusy_320 = {1{1'b0}};
//  assign io_cyclesChannelBusy_321 = {1{1'b0}};
//  assign io_cyclesChannelBusy_322 = {1{1'b0}};
//  assign io_cyclesChannelBusy_323 = {1{1'b0}};
//  assign io_cyclesChannelBusy_324 = {1{1'b0}};
//  assign io_cyclesChannelBusy_325 = {1{1'b0}};
//  assign io_cyclesChannelBusy_326 = {1{1'b0}};
//  assign io_cyclesChannelBusy_327 = {1{1'b0}};
//  assign io_cyclesChannelBusy_328 = {1{1'b0}};
//  assign io_cyclesChannelBusy_329 = {1{1'b0}};
//  assign io_cyclesChannelBusy_330 = {1{1'b0}};
//  assign io_cyclesChannelBusy_331 = {1{1'b0}};
//  assign io_cyclesChannelBusy_332 = {1{1'b0}};
//  assign io_cyclesChannelBusy_333 = {1{1'b0}};
//  assign io_cyclesChannelBusy_334 = {1{1'b0}};
//  assign io_cyclesChannelBusy_335 = {1{1'b0}};
//  assign io_cyclesChannelBusy_336 = {1{1'b0}};
//  assign io_cyclesChannelBusy_337 = {1{1'b0}};
//  assign io_cyclesChannelBusy_338 = {1{1'b0}};
//  assign io_cyclesChannelBusy_339 = {1{1'b0}};
//  assign io_cyclesChannelBusy_340 = {1{1'b0}};
//  assign io_cyclesChannelBusy_341 = {1{1'b0}};
//  assign io_cyclesChannelBusy_342 = {1{1'b0}};
//  assign io_cyclesChannelBusy_343 = {1{1'b0}};
//  assign io_cyclesChannelBusy_344 = {1{1'b0}};
//  assign io_cyclesChannelBusy_345 = {1{1'b0}};
//  assign io_cyclesChannelBusy_346 = {1{1'b0}};
//  assign io_cyclesChannelBusy_347 = {1{1'b0}};
//  assign io_cyclesChannelBusy_348 = {1{1'b0}};
//  assign io_cyclesChannelBusy_349 = {1{1'b0}};
//  assign io_cyclesChannelBusy_350 = {1{1'b0}};
//  assign io_cyclesChannelBusy_351 = {1{1'b0}};
//  assign io_cyclesChannelBusy_352 = {1{1'b0}};
//  assign io_cyclesChannelBusy_353 = {1{1'b0}};
//  assign io_cyclesChannelBusy_354 = {1{1'b0}};
//  assign io_cyclesChannelBusy_355 = {1{1'b0}};
//  assign io_cyclesChannelBusy_356 = {1{1'b0}};
//  assign io_cyclesChannelBusy_357 = {1{1'b0}};
//  assign io_cyclesChannelBusy_358 = {1{1'b0}};
//  assign io_cyclesChannelBusy_359 = {1{1'b0}};
//  assign io_cyclesChannelBusy_360 = {1{1'b0}};
//  assign io_cyclesChannelBusy_361 = {1{1'b0}};
//  assign io_cyclesChannelBusy_362 = {1{1'b0}};
//  assign io_cyclesChannelBusy_363 = {1{1'b0}};
//  assign io_cyclesChannelBusy_364 = {1{1'b0}};
//  assign io_cyclesChannelBusy_365 = {1{1'b0}};
//  assign io_cyclesChannelBusy_366 = {1{1'b0}};
//  assign io_cyclesChannelBusy_367 = {1{1'b0}};
//  assign io_cyclesChannelBusy_368 = {1{1'b0}};
//  assign io_cyclesChannelBusy_369 = {1{1'b0}};
//  assign io_cyclesChannelBusy_370 = {1{1'b0}};
//  assign io_cyclesChannelBusy_371 = {1{1'b0}};
//  assign io_cyclesChannelBusy_372 = {1{1'b0}};
//  assign io_cyclesChannelBusy_373 = {1{1'b0}};
//  assign io_cyclesChannelBusy_374 = {1{1'b0}};
//  assign io_cyclesChannelBusy_375 = {1{1'b0}};
//  assign io_cyclesChannelBusy_376 = {1{1'b0}};
//  assign io_cyclesChannelBusy_377 = {1{1'b0}};
//  assign io_cyclesChannelBusy_378 = {1{1'b0}};
//  assign io_cyclesChannelBusy_379 = {1{1'b0}};
//  assign io_cyclesChannelBusy_380 = {1{1'b0}};
//  assign io_cyclesChannelBusy_381 = {1{1'b0}};
//  assign io_cyclesChannelBusy_382 = {1{1'b0}};
//  assign io_cyclesChannelBusy_383 = {1{1'b0}};
//  assign io_cyclesChannelBusy_384 = {1{1'b0}};
//  assign io_cyclesChannelBusy_385 = {1{1'b0}};
//  assign io_cyclesChannelBusy_386 = {1{1'b0}};
//  assign io_cyclesChannelBusy_387 = {1{1'b0}};
//  assign io_cyclesChannelBusy_388 = {1{1'b0}};
//  assign io_cyclesChannelBusy_389 = {1{1'b0}};
//  assign io_cyclesChannelBusy_390 = {1{1'b0}};
//  assign io_cyclesChannelBusy_391 = {1{1'b0}};
//  assign io_cyclesChannelBusy_392 = {1{1'b0}};
//  assign io_cyclesChannelBusy_393 = {1{1'b0}};
//  assign io_cyclesChannelBusy_394 = {1{1'b0}};
//  assign io_cyclesChannelBusy_395 = {1{1'b0}};
//  assign io_cyclesChannelBusy_396 = {1{1'b0}};
//  assign io_cyclesChannelBusy_397 = {1{1'b0}};
//  assign io_cyclesChannelBusy_398 = {1{1'b0}};
//  assign io_cyclesChannelBusy_399 = {1{1'b0}};
//  assign io_cyclesChannelBusy_400 = {1{1'b0}};
//  assign io_cyclesChannelBusy_401 = {1{1'b0}};
//  assign io_cyclesChannelBusy_402 = {1{1'b0}};
//  assign io_cyclesChannelBusy_403 = {1{1'b0}};
//  assign io_cyclesChannelBusy_404 = {1{1'b0}};
//  assign io_cyclesChannelBusy_405 = {1{1'b0}};
//  assign io_cyclesChannelBusy_406 = {1{1'b0}};
//  assign io_cyclesChannelBusy_407 = {1{1'b0}};
//  assign io_cyclesChannelBusy_408 = {1{1'b0}};
//  assign io_cyclesChannelBusy_409 = {1{1'b0}};
//  assign io_cyclesChannelBusy_410 = {1{1'b0}};
//  assign io_cyclesChannelBusy_411 = {1{1'b0}};
//  assign io_cyclesChannelBusy_412 = {1{1'b0}};
//  assign io_cyclesChannelBusy_413 = {1{1'b0}};
//  assign io_cyclesChannelBusy_414 = {1{1'b0}};
//  assign io_cyclesChannelBusy_415 = {1{1'b0}};
//  assign io_cyclesChannelBusy_416 = {1{1'b0}};
//  assign io_cyclesChannelBusy_417 = {1{1'b0}};
//  assign io_cyclesChannelBusy_418 = {1{1'b0}};
//  assign io_cyclesChannelBusy_419 = {1{1'b0}};
//  assign io_cyclesChannelBusy_420 = {1{1'b0}};
//  assign io_cyclesChannelBusy_421 = {1{1'b0}};
//  assign io_cyclesChannelBusy_422 = {1{1'b0}};
//  assign io_cyclesChannelBusy_423 = {1{1'b0}};
//  assign io_cyclesChannelBusy_424 = {1{1'b0}};
//  assign io_cyclesChannelBusy_425 = {1{1'b0}};
//  assign io_cyclesChannelBusy_426 = {1{1'b0}};
//  assign io_cyclesChannelBusy_427 = {1{1'b0}};
//  assign io_cyclesChannelBusy_428 = {1{1'b0}};
//  assign io_cyclesChannelBusy_429 = {1{1'b0}};
//  assign io_cyclesChannelBusy_430 = {1{1'b0}};
//  assign io_cyclesChannelBusy_431 = {1{1'b0}};
//  assign io_cyclesChannelBusy_432 = {1{1'b0}};
//  assign io_cyclesChannelBusy_433 = {1{1'b0}};
//  assign io_cyclesChannelBusy_434 = {1{1'b0}};
//  assign io_cyclesChannelBusy_435 = {1{1'b0}};
//  assign io_cyclesChannelBusy_436 = {1{1'b0}};
//  assign io_cyclesChannelBusy_437 = {1{1'b0}};
//  assign io_cyclesChannelBusy_438 = {1{1'b0}};
//  assign io_cyclesChannelBusy_439 = {1{1'b0}};
//  assign io_cyclesChannelBusy_440 = {1{1'b0}};
//  assign io_cyclesChannelBusy_441 = {1{1'b0}};
//  assign io_cyclesChannelBusy_442 = {1{1'b0}};
//  assign io_cyclesChannelBusy_443 = {1{1'b0}};
//  assign io_cyclesChannelBusy_444 = {1{1'b0}};
//  assign io_cyclesChannelBusy_445 = {1{1'b0}};
//  assign io_cyclesChannelBusy_446 = {1{1'b0}};
//  assign io_cyclesChannelBusy_447 = {1{1'b0}};
//  assign io_cyclesChannelBusy_448 = {1{1'b0}};
//  assign io_cyclesChannelBusy_449 = {1{1'b0}};
//  assign io_cyclesChannelBusy_450 = {1{1'b0}};
//  assign io_cyclesChannelBusy_451 = {1{1'b0}};
//  assign io_cyclesChannelBusy_452 = {1{1'b0}};
//  assign io_cyclesChannelBusy_453 = {1{1'b0}};
//  assign io_cyclesChannelBusy_454 = {1{1'b0}};
//  assign io_cyclesChannelBusy_455 = {1{1'b0}};
//  assign io_cyclesChannelBusy_456 = {1{1'b0}};
//  assign io_cyclesChannelBusy_457 = {1{1'b0}};
//  assign io_cyclesChannelBusy_458 = {1{1'b0}};
//  assign io_cyclesChannelBusy_459 = {1{1'b0}};
//  assign io_cyclesChannelBusy_460 = {1{1'b0}};
//  assign io_cyclesChannelBusy_461 = {1{1'b0}};
//  assign io_cyclesChannelBusy_462 = {1{1'b0}};
//  assign io_cyclesChannelBusy_463 = {1{1'b0}};
//  assign io_cyclesChannelBusy_464 = {1{1'b0}};
//  assign io_cyclesChannelBusy_465 = {1{1'b0}};
//  assign io_cyclesChannelBusy_466 = {1{1'b0}};
//  assign io_cyclesChannelBusy_467 = {1{1'b0}};
//  assign io_cyclesChannelBusy_468 = {1{1'b0}};
//  assign io_cyclesChannelBusy_469 = {1{1'b0}};
//  assign io_cyclesChannelBusy_470 = {1{1'b0}};
//  assign io_cyclesChannelBusy_471 = {1{1'b0}};
//  assign io_cyclesChannelBusy_472 = {1{1'b0}};
//  assign io_cyclesChannelBusy_473 = {1{1'b0}};
//  assign io_cyclesChannelBusy_474 = {1{1'b0}};
//  assign io_cyclesChannelBusy_475 = {1{1'b0}};
//  assign io_cyclesChannelBusy_476 = {1{1'b0}};
//  assign io_cyclesChannelBusy_477 = {1{1'b0}};
//  assign io_cyclesChannelBusy_478 = {1{1'b0}};
//  assign io_cyclesChannelBusy_479 = {1{1'b0}};
//  assign io_cyclesChannelBusy_480 = {1{1'b0}};
//  assign io_cyclesChannelBusy_481 = {1{1'b0}};
//  assign io_cyclesChannelBusy_482 = {1{1'b0}};
//  assign io_cyclesChannelBusy_483 = {1{1'b0}};
//  assign io_cyclesChannelBusy_484 = {1{1'b0}};
//  assign io_cyclesChannelBusy_485 = {1{1'b0}};
//  assign io_cyclesChannelBusy_486 = {1{1'b0}};
//  assign io_cyclesChannelBusy_487 = {1{1'b0}};
//  assign io_cyclesChannelBusy_488 = {1{1'b0}};
//  assign io_cyclesChannelBusy_489 = {1{1'b0}};
//  assign io_cyclesChannelBusy_490 = {1{1'b0}};
//  assign io_cyclesChannelBusy_491 = {1{1'b0}};
//  assign io_cyclesChannelBusy_492 = {1{1'b0}};
//  assign io_cyclesChannelBusy_493 = {1{1'b0}};
//  assign io_cyclesChannelBusy_494 = {1{1'b0}};
//  assign io_cyclesChannelBusy_495 = {1{1'b0}};
//  assign io_cyclesChannelBusy_496 = {1{1'b0}};
//  assign io_cyclesChannelBusy_497 = {1{1'b0}};
//  assign io_cyclesChannelBusy_498 = {1{1'b0}};
//  assign io_cyclesChannelBusy_499 = {1{1'b0}};
//  assign io_cyclesChannelBusy_500 = {1{1'b0}};
//  assign io_cyclesChannelBusy_501 = {1{1'b0}};
//  assign io_cyclesChannelBusy_502 = {1{1'b0}};
//  assign io_cyclesChannelBusy_503 = {1{1'b0}};
//  assign io_cyclesChannelBusy_504 = {1{1'b0}};
//  assign io_cyclesChannelBusy_505 = {1{1'b0}};
//  assign io_cyclesChannelBusy_506 = {1{1'b0}};
//  assign io_cyclesChannelBusy_507 = {1{1'b0}};
//  assign io_cyclesChannelBusy_508 = {1{1'b0}};
//  assign io_cyclesChannelBusy_509 = {1{1'b0}};
//  assign io_cyclesChannelBusy_510 = {1{1'b0}};
//  assign io_cyclesChannelBusy_511 = {1{1'b0}};
//  assign io_cyclesChannelBusy_512 = {1{1'b0}};
//  assign io_cyclesChannelBusy_513 = {1{1'b0}};
//  assign io_cyclesChannelBusy_514 = {1{1'b0}};
//  assign io_cyclesChannelBusy_515 = {1{1'b0}};
//  assign io_cyclesChannelBusy_516 = {1{1'b0}};
//  assign io_cyclesChannelBusy_517 = {1{1'b0}};
//  assign io_cyclesChannelBusy_518 = {1{1'b0}};
//  assign io_cyclesChannelBusy_519 = {1{1'b0}};
//  assign io_cyclesChannelBusy_520 = {1{1'b0}};
//  assign io_cyclesChannelBusy_521 = {1{1'b0}};
//  assign io_cyclesChannelBusy_522 = {1{1'b0}};
//  assign io_cyclesChannelBusy_523 = {1{1'b0}};
//  assign io_cyclesChannelBusy_524 = {1{1'b0}};
//  assign io_cyclesChannelBusy_525 = {1{1'b0}};
//  assign io_cyclesChannelBusy_526 = {1{1'b0}};
//  assign io_cyclesChannelBusy_527 = {1{1'b0}};
//  assign io_cyclesChannelBusy_528 = {1{1'b0}};
//  assign io_cyclesChannelBusy_529 = {1{1'b0}};
//  assign io_cyclesChannelBusy_530 = {1{1'b0}};
//  assign io_cyclesChannelBusy_531 = {1{1'b0}};
//  assign io_cyclesChannelBusy_532 = {1{1'b0}};
//  assign io_cyclesChannelBusy_533 = {1{1'b0}};
//  assign io_cyclesChannelBusy_534 = {1{1'b0}};
//  assign io_cyclesChannelBusy_535 = {1{1'b0}};
//  assign io_cyclesChannelBusy_536 = {1{1'b0}};
//  assign io_cyclesChannelBusy_537 = {1{1'b0}};
//  assign io_cyclesChannelBusy_538 = {1{1'b0}};
//  assign io_cyclesChannelBusy_539 = {1{1'b0}};
//  assign io_cyclesChannelBusy_540 = {1{1'b0}};
//  assign io_cyclesChannelBusy_541 = {1{1'b0}};
//  assign io_cyclesChannelBusy_542 = {1{1'b0}};
//  assign io_cyclesChannelBusy_543 = {1{1'b0}};
//  assign io_cyclesChannelBusy_544 = {1{1'b0}};
//  assign io_cyclesChannelBusy_545 = {1{1'b0}};
//  assign io_cyclesChannelBusy_546 = {1{1'b0}};
//  assign io_cyclesChannelBusy_547 = {1{1'b0}};
//  assign io_cyclesChannelBusy_548 = {1{1'b0}};
//  assign io_cyclesChannelBusy_549 = {1{1'b0}};
//  assign io_cyclesChannelBusy_550 = {1{1'b0}};
//  assign io_cyclesChannelBusy_551 = {1{1'b0}};
//  assign io_cyclesChannelBusy_552 = {1{1'b0}};
//  assign io_cyclesChannelBusy_553 = {1{1'b0}};
//  assign io_cyclesChannelBusy_554 = {1{1'b0}};
//  assign io_cyclesChannelBusy_555 = {1{1'b0}};
//  assign io_cyclesChannelBusy_556 = {1{1'b0}};
//  assign io_cyclesChannelBusy_557 = {1{1'b0}};
//  assign io_cyclesChannelBusy_558 = {1{1'b0}};
//  assign io_cyclesChannelBusy_559 = {1{1'b0}};
//  assign io_cyclesChannelBusy_560 = {1{1'b0}};
//  assign io_cyclesChannelBusy_561 = {1{1'b0}};
//  assign io_cyclesChannelBusy_562 = {1{1'b0}};
//  assign io_cyclesChannelBusy_563 = {1{1'b0}};
//  assign io_cyclesChannelBusy_564 = {1{1'b0}};
//  assign io_cyclesChannelBusy_565 = {1{1'b0}};
//  assign io_cyclesChannelBusy_566 = {1{1'b0}};
//  assign io_cyclesChannelBusy_567 = {1{1'b0}};
//  assign io_cyclesChannelBusy_568 = {1{1'b0}};
//  assign io_cyclesChannelBusy_569 = {1{1'b0}};
//  assign io_cyclesChannelBusy_570 = {1{1'b0}};
//  assign io_cyclesChannelBusy_571 = {1{1'b0}};
//  assign io_cyclesChannelBusy_572 = {1{1'b0}};
//  assign io_cyclesChannelBusy_573 = {1{1'b0}};
//  assign io_cyclesChannelBusy_574 = {1{1'b0}};
//  assign io_cyclesChannelBusy_575 = {1{1'b0}};
//  assign io_cyclesChannelBusy_576 = {1{1'b0}};
//  assign io_cyclesChannelBusy_577 = {1{1'b0}};
//  assign io_cyclesChannelBusy_578 = {1{1'b0}};
//  assign io_cyclesChannelBusy_579 = {1{1'b0}};
//  assign io_cyclesChannelBusy_580 = {1{1'b0}};
//  assign io_cyclesChannelBusy_581 = {1{1'b0}};
//  assign io_cyclesChannelBusy_582 = {1{1'b0}};
//  assign io_cyclesChannelBusy_583 = {1{1'b0}};
//  assign io_cyclesChannelBusy_584 = {1{1'b0}};
//  assign io_cyclesChannelBusy_585 = {1{1'b0}};
//  assign io_cyclesChannelBusy_586 = {1{1'b0}};
//  assign io_cyclesChannelBusy_587 = {1{1'b0}};
//  assign io_cyclesChannelBusy_588 = {1{1'b0}};
//  assign io_cyclesChannelBusy_589 = {1{1'b0}};
//  assign io_cyclesChannelBusy_590 = {1{1'b0}};
//  assign io_cyclesChannelBusy_591 = {1{1'b0}};
//  assign io_cyclesChannelBusy_592 = {1{1'b0}};
//  assign io_cyclesChannelBusy_593 = {1{1'b0}};
//  assign io_cyclesChannelBusy_594 = {1{1'b0}};
//  assign io_cyclesChannelBusy_595 = {1{1'b0}};
//  assign io_cyclesChannelBusy_596 = {1{1'b0}};
//  assign io_cyclesChannelBusy_597 = {1{1'b0}};
//  assign io_cyclesChannelBusy_598 = {1{1'b0}};
//  assign io_cyclesChannelBusy_599 = {1{1'b0}};
//  assign io_cyclesChannelBusy_600 = {1{1'b0}};
//  assign io_cyclesChannelBusy_601 = {1{1'b0}};
//  assign io_cyclesChannelBusy_602 = {1{1'b0}};
//  assign io_cyclesChannelBusy_603 = {1{1'b0}};
//  assign io_cyclesChannelBusy_604 = {1{1'b0}};
//  assign io_cyclesChannelBusy_605 = {1{1'b0}};
//  assign io_cyclesChannelBusy_606 = {1{1'b0}};
//  assign io_cyclesChannelBusy_607 = {1{1'b0}};
//  assign io_cyclesChannelBusy_608 = {1{1'b0}};
//  assign io_cyclesChannelBusy_609 = {1{1'b0}};
//  assign io_cyclesChannelBusy_610 = {1{1'b0}};
//  assign io_cyclesChannelBusy_611 = {1{1'b0}};
//  assign io_cyclesChannelBusy_612 = {1{1'b0}};
//  assign io_cyclesChannelBusy_613 = {1{1'b0}};
//  assign io_cyclesChannelBusy_614 = {1{1'b0}};
//  assign io_cyclesChannelBusy_615 = {1{1'b0}};
//  assign io_cyclesChannelBusy_616 = {1{1'b0}};
//  assign io_cyclesChannelBusy_617 = {1{1'b0}};
//  assign io_cyclesChannelBusy_618 = {1{1'b0}};
//  assign io_cyclesChannelBusy_619 = {1{1'b0}};
//  assign io_cyclesChannelBusy_620 = {1{1'b0}};
//  assign io_cyclesChannelBusy_621 = {1{1'b0}};
//  assign io_cyclesChannelBusy_622 = {1{1'b0}};
//  assign io_cyclesChannelBusy_623 = {1{1'b0}};
//  assign io_cyclesChannelBusy_624 = {1{1'b0}};
//  assign io_cyclesChannelBusy_625 = {1{1'b0}};
//  assign io_cyclesChannelBusy_626 = {1{1'b0}};
//  assign io_cyclesChannelBusy_627 = {1{1'b0}};
//  assign io_cyclesChannelBusy_628 = {1{1'b0}};
//  assign io_cyclesChannelBusy_629 = {1{1'b0}};
//  assign io_cyclesChannelBusy_630 = {1{1'b0}};
//  assign io_cyclesChannelBusy_631 = {1{1'b0}};
//  assign io_cyclesChannelBusy_632 = {1{1'b0}};
//  assign io_cyclesChannelBusy_633 = {1{1'b0}};
//  assign io_cyclesChannelBusy_634 = {1{1'b0}};
//  assign io_cyclesChannelBusy_635 = {1{1'b0}};
//  assign io_cyclesChannelBusy_636 = {1{1'b0}};
//  assign io_cyclesChannelBusy_637 = {1{1'b0}};
//  assign io_cyclesChannelBusy_638 = {1{1'b0}};
//  assign io_cyclesChannelBusy_639 = {1{1'b0}};
//  assign io_cyclesRouterBusy_3 = {1{1'b0}};
//  assign io_cyclesRouterBusy_4 = {1{1'b0}};
//  assign io_cyclesRouterBusy_5 = {1{1'b0}};
//  assign io_cyclesRouterBusy_6 = {1{1'b0}};
//  assign io_cyclesRouterBusy_7 = {1{1'b0}};
//  assign io_cyclesRouterBusy_8 = {1{1'b0}};
//  assign io_cyclesRouterBusy_9 = {1{1'b0}};
//  assign io_cyclesRouterBusy_10 = {1{1'b0}};
//  assign io_cyclesRouterBusy_11 = {1{1'b0}};
//  assign io_cyclesRouterBusy_12 = {1{1'b0}};
//  assign io_cyclesRouterBusy_13 = {1{1'b0}};
//  assign io_cyclesRouterBusy_14 = {1{1'b0}};
//  assign io_cyclesRouterBusy_15 = {1{1'b0}};
//  assign io_cyclesRouterBusy_16 = {1{1'b0}};
//  assign io_cyclesRouterBusy_17 = {1{1'b0}};
//  assign io_cyclesRouterBusy_18 = {1{1'b0}};
//  assign io_cyclesRouterBusy_19 = {1{1'b0}};
//  assign io_cyclesRouterBusy_20 = {1{1'b0}};
//  assign io_cyclesRouterBusy_21 = {1{1'b0}};
//  assign io_cyclesRouterBusy_22 = {1{1'b0}};
//  assign io_cyclesRouterBusy_23 = {1{1'b0}};
//  assign io_cyclesRouterBusy_24 = {1{1'b0}};
//  assign io_cyclesRouterBusy_25 = {1{1'b0}};
//  assign io_cyclesRouterBusy_26 = {1{1'b0}};
//  assign io_cyclesRouterBusy_27 = {1{1'b0}};
//  assign io_cyclesRouterBusy_28 = {1{1'b0}};
//  assign io_cyclesRouterBusy_29 = {1{1'b0}};
//  assign io_cyclesRouterBusy_30 = {1{1'b0}};
//  assign io_cyclesRouterBusy_31 = {1{1'b0}};
//  assign io_cyclesRouterBusy_32 = {1{1'b0}};
//  assign io_cyclesRouterBusy_33 = {1{1'b0}};
//  assign io_cyclesRouterBusy_34 = {1{1'b0}};
//  assign io_cyclesRouterBusy_35 = {1{1'b0}};
//  assign io_cyclesRouterBusy_36 = {1{1'b0}};
//  assign io_cyclesRouterBusy_37 = {1{1'b0}};
//  assign io_cyclesRouterBusy_38 = {1{1'b0}};
//  assign io_cyclesRouterBusy_39 = {1{1'b0}};
//  assign io_cyclesRouterBusy_40 = {1{1'b0}};
//  assign io_cyclesRouterBusy_41 = {1{1'b0}};
//  assign io_cyclesRouterBusy_42 = {1{1'b0}};
//  assign io_cyclesRouterBusy_43 = {1{1'b0}};
//  assign io_cyclesRouterBusy_44 = {1{1'b0}};
//  assign io_cyclesRouterBusy_45 = {1{1'b0}};
//  assign io_cyclesRouterBusy_46 = {1{1'b0}};
//  assign io_cyclesRouterBusy_47 = {1{1'b0}};
//  assign io_cyclesRouterBusy_48 = {1{1'b0}};
//  assign io_cyclesRouterBusy_49 = {1{1'b0}};
//  assign io_cyclesRouterBusy_50 = {1{1'b0}};
//  assign io_cyclesRouterBusy_51 = {1{1'b0}};
//  assign io_cyclesRouterBusy_52 = {1{1'b0}};
//  assign io_cyclesRouterBusy_53 = {1{1'b0}};
//  assign io_cyclesRouterBusy_54 = {1{1'b0}};
//  assign io_cyclesRouterBusy_55 = {1{1'b0}};
//  assign io_cyclesRouterBusy_56 = {1{1'b0}};
//  assign io_cyclesRouterBusy_57 = {1{1'b0}};
//  assign io_cyclesRouterBusy_58 = {1{1'b0}};
//  assign io_cyclesRouterBusy_59 = {1{1'b0}};
//  assign io_cyclesRouterBusy_60 = {1{1'b0}};
//  assign io_cyclesRouterBusy_61 = {1{1'b0}};
//  assign io_cyclesRouterBusy_62 = {1{1'b0}};
//  assign io_cyclesRouterBusy_63 = {1{1'b0}};
//  assign io_cyclesRouterBusy_64 = {1{1'b0}};
//  assign io_cyclesRouterBusy_65 = {1{1'b0}};
//  assign io_cyclesRouterBusy_66 = {1{1'b0}};
//  assign io_cyclesRouterBusy_67 = {1{1'b0}};
//  assign io_cyclesRouterBusy_68 = {1{1'b0}};
//  assign io_cyclesRouterBusy_69 = {1{1'b0}};
//  assign io_cyclesRouterBusy_70 = {1{1'b0}};
//  assign io_cyclesRouterBusy_71 = {1{1'b0}};
//  assign io_cyclesRouterBusy_72 = {1{1'b0}};
//  assign io_cyclesRouterBusy_73 = {1{1'b0}};
//  assign io_cyclesRouterBusy_74 = {1{1'b0}};
//  assign io_cyclesRouterBusy_75 = {1{1'b0}};
//  assign io_cyclesRouterBusy_76 = {1{1'b0}};
//  assign io_cyclesRouterBusy_77 = {1{1'b0}};
//  assign io_cyclesRouterBusy_78 = {1{1'b0}};
//  assign io_cyclesRouterBusy_79 = {1{1'b0}};
//  assign io_cyclesRouterBusy_80 = {1{1'b0}};
//  assign io_cyclesRouterBusy_81 = {1{1'b0}};
//  assign io_cyclesRouterBusy_82 = {1{1'b0}};
//  assign io_cyclesRouterBusy_83 = {1{1'b0}};
//  assign io_cyclesRouterBusy_84 = {1{1'b0}};
//  assign io_cyclesRouterBusy_85 = {1{1'b0}};
//  assign io_cyclesRouterBusy_86 = {1{1'b0}};
//  assign io_cyclesRouterBusy_87 = {1{1'b0}};
//  assign io_cyclesRouterBusy_88 = {1{1'b0}};
//  assign io_cyclesRouterBusy_89 = {1{1'b0}};
//  assign io_cyclesRouterBusy_90 = {1{1'b0}};
//  assign io_cyclesRouterBusy_91 = {1{1'b0}};
//  assign io_cyclesRouterBusy_92 = {1{1'b0}};
//  assign io_cyclesRouterBusy_93 = {1{1'b0}};
//  assign io_cyclesRouterBusy_94 = {1{1'b0}};
//  assign io_cyclesRouterBusy_95 = {1{1'b0}};
//  assign io_cyclesRouterBusy_96 = {1{1'b0}};
//  assign io_cyclesRouterBusy_97 = {1{1'b0}};
//  assign io_cyclesRouterBusy_98 = {1{1'b0}};
//  assign io_cyclesRouterBusy_99 = {1{1'b0}};
//  assign io_cyclesRouterBusy_100 = {1{1'b0}};
//  assign io_cyclesRouterBusy_101 = {1{1'b0}};
//  assign io_cyclesRouterBusy_102 = {1{1'b0}};
//  assign io_cyclesRouterBusy_103 = {1{1'b0}};
//  assign io_cyclesRouterBusy_104 = {1{1'b0}};
//  assign io_cyclesRouterBusy_105 = {1{1'b0}};
//  assign io_cyclesRouterBusy_106 = {1{1'b0}};
//  assign io_cyclesRouterBusy_107 = {1{1'b0}};
//  assign io_cyclesRouterBusy_108 = {1{1'b0}};
//  assign io_cyclesRouterBusy_109 = {1{1'b0}};
//  assign io_cyclesRouterBusy_110 = {1{1'b0}};
//  assign io_cyclesRouterBusy_111 = {1{1'b0}};
//  assign io_cyclesRouterBusy_112 = {1{1'b0}};
//  assign io_cyclesRouterBusy_113 = {1{1'b0}};
//  assign io_cyclesRouterBusy_114 = {1{1'b0}};
//  assign io_cyclesRouterBusy_115 = {1{1'b0}};
//  assign io_cyclesRouterBusy_116 = {1{1'b0}};
//  assign io_cyclesRouterBusy_117 = {1{1'b0}};
//  assign io_cyclesRouterBusy_118 = {1{1'b0}};
//  assign io_cyclesRouterBusy_119 = {1{1'b0}};
//  assign io_cyclesRouterBusy_120 = {1{1'b0}};
//  assign io_cyclesRouterBusy_121 = {1{1'b0}};
//  assign io_cyclesRouterBusy_122 = {1{1'b0}};
//  assign io_cyclesRouterBusy_123 = {1{1'b0}};
//  assign io_cyclesRouterBusy_124 = {1{1'b0}};
//  assign io_cyclesRouterBusy_125 = {1{1'b0}};
//  assign io_cyclesRouterBusy_126 = {1{1'b0}};
//  assign io_cyclesRouterBusy_127 = {1{1'b0}};
// synthesis translate_on
`endif
  assign io_cyclesChannelBusy_1 = BusProbe_io_cyclesChannelBusy_1;
  assign io_cyclesChannelBusy_6 = BusProbe_1_io_cyclesChannelBusy_1;
  assign io_cyclesChannelBusy_7 = BusProbe_1_io_cyclesChannelBusy_2;
  assign io_cyclesChannelBusy_12 = BusProbe_2_io_cyclesChannelBusy_2;
  assign io_cyclesRouterBusy_0 = BusProbe_1_io_cyclesRouterBusy;
  assign io_cyclesRouterBusy_1 = BusProbe_2_io_cyclesRouterBusy;
  assign io_cyclesRouterBusy_2 = BusProbe_io_cyclesRouterBusy;
  assign io_outChannels_0_flitValid = VCRouterWrapper_io_outChannels_0_flitValid;
  assign io_outChannels_0_flit_x = VCRouterWrapper_io_outChannels_0_flit_x;
  assign io_outChannels_1_flitValid = VCRouterWrapper_1_io_outChannels_0_flitValid;
  assign io_outChannels_1_flit_x = VCRouterWrapper_1_io_outChannels_0_flit_x;
  assign io_outChannels_2_flitValid = VCRouterWrapper_2_io_outChannels_0_flitValid;
  assign io_outChannels_2_flit_x = VCRouterWrapper_2_io_outChannels_0_flit_x;
  assign io_inChannels_0_credit_0_grant = VCRouterWrapper_io_inChannels_0_credit_0_grant;
  assign io_inChannels_0_credit_1_grant = VCRouterWrapper_io_inChannels_0_credit_1_grant;
  assign io_inChannels_1_credit_0_grant = VCRouterWrapper_1_io_inChannels_0_credit_0_grant;
  assign io_inChannels_1_credit_1_grant = VCRouterWrapper_1_io_inChannels_0_credit_1_grant;
  assign io_inChannels_2_credit_0_grant = VCRouterWrapper_2_io_inChannels_0_credit_0_grant;
  assign io_inChannels_2_credit_1_grant = VCRouterWrapper_2_io_inChannels_0_credit_1_grant;
  VCRouterWrapper_0 VCRouterWrapper(.clk(clk), .reset(reset),
       .io_inChannels_4_flit_x( OpenSoC_VCConstantEndpoint_2_io_outChannels_4_flit_x ),
       .io_inChannels_4_flitValid( OpenSoC_VCConstantEndpoint_2_io_outChannels_4_flitValid ),
       .io_inChannels_4_credit_1_grant( VCRouterWrapper_io_inChannels_4_credit_1_grant ),
       .io_inChannels_4_credit_0_grant( VCRouterWrapper_io_inChannels_4_credit_0_grant ),
       .io_inChannels_3_flit_x( OpenSoC_VCConstantEndpoint_1_io_outChannels_3_flit_x ),
       .io_inChannels_3_flitValid( OpenSoC_VCConstantEndpoint_1_io_outChannels_3_flitValid ),
       .io_inChannels_3_credit_1_grant( VCRouterWrapper_io_inChannels_3_credit_1_grant ),
       .io_inChannels_3_credit_0_grant( VCRouterWrapper_io_inChannels_3_credit_0_grant ),
       .io_inChannels_2_flit_x( CreditBuffer_1_io_out_2_flit_x ),
       .io_inChannels_2_flitValid( CreditBuffer_1_io_out_2_flitValid ),
       .io_inChannels_2_credit_1_grant( VCRouterWrapper_io_inChannels_2_credit_1_grant ),
       .io_inChannels_2_credit_0_grant( VCRouterWrapper_io_inChannels_2_credit_0_grant ),
       .io_inChannels_1_flit_x( OpenSoC_VCConstantEndpoint_io_outChannels_1_flit_x ),
       .io_inChannels_1_flitValid( OpenSoC_VCConstantEndpoint_io_outChannels_1_flitValid ),
       .io_inChannels_1_credit_1_grant( VCRouterWrapper_io_inChannels_1_credit_1_grant ),
       .io_inChannels_1_credit_0_grant( VCRouterWrapper_io_inChannels_1_credit_0_grant ),
       .io_inChannels_0_flit_x( io_inChannels_0_flit_x ),
       .io_inChannels_0_flitValid( io_inChannels_0_flitValid ),
       .io_inChannels_0_credit_1_grant( VCRouterWrapper_io_inChannels_0_credit_1_grant ),
       .io_inChannels_0_credit_0_grant( VCRouterWrapper_io_inChannels_0_credit_0_grant ),
       .io_outChannels_4_flit_x( VCRouterWrapper_io_outChannels_4_flit_x ),
       .io_outChannels_4_flitValid( VCRouterWrapper_io_outChannels_4_flitValid ),
       //.io_outChannels_4_credit_1_grant(  )
       //.io_outChannels_4_credit_0_grant(  )
       .io_outChannels_3_flit_x( VCRouterWrapper_io_outChannels_3_flit_x ),
       .io_outChannels_3_flitValid( VCRouterWrapper_io_outChannels_3_flitValid ),
       //.io_outChannels_3_credit_1_grant(  )
       //.io_outChannels_3_credit_0_grant(  )
       //.io_outChannels_2_flit_x(  )
       //.io_outChannels_2_flitValid(  )
       //.io_outChannels_2_credit_1_grant(  )
       //.io_outChannels_2_credit_0_grant(  )
       .io_outChannels_1_flit_x( VCRouterWrapper_io_outChannels_1_flit_x ),
       .io_outChannels_1_flitValid( VCRouterWrapper_io_outChannels_1_flitValid ),
       .io_outChannels_1_credit_1_grant( CreditBuffer_io_in_1_credit_1_grant ),
       .io_outChannels_1_credit_0_grant( CreditBuffer_io_in_1_credit_0_grant ),
       .io_outChannels_0_flit_x( VCRouterWrapper_io_outChannels_0_flit_x ),
       .io_outChannels_0_flitValid( VCRouterWrapper_io_outChannels_0_flitValid ),
       .io_outChannels_0_credit_1_grant( io_outChannels_0_credit_1_grant ),
       .io_outChannels_0_credit_0_grant( io_outChannels_0_credit_0_grant ),
       //.io_counters_1_counterVal(  )
       //.io_counters_1_counterIndex(  )
       //.io_counters_0_counterVal(  )
       //.io_counters_0_counterIndex(  )
       .io_bypass( io_bypass_0 )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign VCRouterWrapper.io_outChannels_4_credit_1_grant = {1{1'b0}};
    assign VCRouterWrapper.io_outChannels_4_credit_0_grant = {1{1'b0}};
    assign VCRouterWrapper.io_outChannels_3_credit_1_grant = {1{1'b0}};
    assign VCRouterWrapper.io_outChannels_3_credit_0_grant = {1{1'b0}};
    assign VCRouterWrapper.io_outChannels_2_credit_1_grant = {1{1'b0}};
    assign VCRouterWrapper.io_outChannels_2_credit_0_grant = {1{1'b0}};
// synthesis translate_on
`endif
  BusProbe_0 BusProbe(.clk(clk), .reset(reset),
       //.io_inFlit_4_x(  )
       //.io_inFlit_3_x(  )
       //.io_inFlit_2_x(  )
       .io_inFlit_1_x( VCRouterWrapper_io_outChannels_1_flit_x ),
       //.io_inFlit_0_x(  )
       //.io_inValid_4(  )
       //.io_inValid_3(  )
       //.io_inValid_2(  )
       .io_inValid_1( VCRouterWrapper_io_outChannels_1_flitValid ),
       //.io_inValid_0(  )
       .io_routerCord( 1'h0 ),
       //.io_startRecording(  )
       //.io_cyclesChannelBusy_4(  )
       //.io_cyclesChannelBusy_3(  )
       //.io_cyclesChannelBusy_2(  )
       .io_cyclesChannelBusy_1( BusProbe_io_cyclesChannelBusy_1 ),
       //.io_cyclesChannelBusy_0(  )
       .io_cyclesRouterBusy( BusProbe_io_cyclesRouterBusy )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign BusProbe.io_inValid_4 = {1{1'b0}};
    assign BusProbe.io_inValid_3 = {1{1'b0}};
    assign BusProbe.io_inValid_2 = {1{1'b0}};
    assign BusProbe.io_inValid_0 = {1{1'b0}};
// synthesis translate_on
`endif
  CreditBuffer CreditBuffer(.clk(clk), .reset(reset),
       //.io_in_4_flit_x(  )
       //.io_in_4_flitValid(  )
       //.io_in_4_credit_1_grant(  )
       //.io_in_4_credit_0_grant(  )
       //.io_in_3_flit_x(  )
       //.io_in_3_flitValid(  )
       //.io_in_3_credit_1_grant(  )
       //.io_in_3_credit_0_grant(  )
       //.io_in_2_flit_x(  )
       //.io_in_2_flitValid(  )
       //.io_in_2_credit_1_grant(  )
       //.io_in_2_credit_0_grant(  )
       .io_in_1_flit_x( VCRouterWrapper_io_outChannels_1_flit_x ),
       .io_in_1_flitValid( VCRouterWrapper_io_outChannels_1_flitValid ),
       .io_in_1_credit_1_grant( CreditBuffer_io_in_1_credit_1_grant ),
       .io_in_1_credit_0_grant( CreditBuffer_io_in_1_credit_0_grant ),
       //.io_in_0_flit_x(  )
       //.io_in_0_flitValid(  )
       //.io_in_0_credit_1_grant(  )
       //.io_in_0_credit_0_grant(  )
       //.io_out_4_flit_x(  )
       //.io_out_4_flitValid(  )
       //.io_out_4_credit_1_grant(  )
       //.io_out_4_credit_0_grant(  )
       //.io_out_3_flit_x(  )
       //.io_out_3_flitValid(  )
       //.io_out_3_credit_1_grant(  )
       //.io_out_3_credit_0_grant(  )
       //.io_out_2_flit_x(  )
       //.io_out_2_flitValid(  )
       //.io_out_2_credit_1_grant(  )
       //.io_out_2_credit_0_grant(  )
       .io_out_1_flit_x( CreditBuffer_io_out_1_flit_x ),
       .io_out_1_flitValid( CreditBuffer_io_out_1_flitValid ),
       .io_out_1_credit_1_grant( VCRouterWrapper_1_io_inChannels_1_credit_1_grant ),
       .io_out_1_credit_0_grant( VCRouterWrapper_1_io_inChannels_1_credit_0_grant )
       //.io_out_0_flit_x(  )
       //.io_out_0_flitValid(  )
       //.io_out_0_credit_1_grant(  )
       //.io_out_0_credit_0_grant(  )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign CreditBuffer.io_in_4_flit_x = {2{1'b0}};
    assign CreditBuffer.io_in_4_flitValid = {1{1'b0}};
    assign CreditBuffer.io_in_3_flit_x = {2{1'b0}};
    assign CreditBuffer.io_in_3_flitValid = {1{1'b0}};
    assign CreditBuffer.io_in_2_flit_x = {2{1'b0}};
    assign CreditBuffer.io_in_2_flitValid = {1{1'b0}};
    assign CreditBuffer.io_in_0_flit_x = {2{1'b0}};
    assign CreditBuffer.io_in_0_flitValid = {1{1'b0}};
    assign CreditBuffer.io_out_4_credit_1_grant = {1{1'b0}};
    assign CreditBuffer.io_out_4_credit_0_grant = {1{1'b0}};
    assign CreditBuffer.io_out_3_credit_1_grant = {1{1'b0}};
    assign CreditBuffer.io_out_3_credit_0_grant = {1{1'b0}};
    assign CreditBuffer.io_out_2_credit_1_grant = {1{1'b0}};
    assign CreditBuffer.io_out_2_credit_0_grant = {1{1'b0}};
    assign CreditBuffer.io_out_0_credit_1_grant = {1{1'b0}};
    assign CreditBuffer.io_out_0_credit_0_grant = {1{1'b0}};
// synthesis translate_on
`endif
  VCRouterWrapper_1 VCRouterWrapper_1(.clk(clk), .reset(reset),
       .io_inChannels_4_flit_x( OpenSoC_VCConstantEndpoint_4_io_outChannels_4_flit_x ),
       .io_inChannels_4_flitValid( OpenSoC_VCConstantEndpoint_4_io_outChannels_4_flitValid ),
       .io_inChannels_4_credit_1_grant( VCRouterWrapper_1_io_inChannels_4_credit_1_grant ),
       .io_inChannels_4_credit_0_grant( VCRouterWrapper_1_io_inChannels_4_credit_0_grant ),
       .io_inChannels_3_flit_x( OpenSoC_VCConstantEndpoint_3_io_outChannels_3_flit_x ),
       .io_inChannels_3_flitValid( OpenSoC_VCConstantEndpoint_3_io_outChannels_3_flitValid ),
       .io_inChannels_3_credit_1_grant( VCRouterWrapper_1_io_inChannels_3_credit_1_grant ),
       .io_inChannels_3_credit_0_grant( VCRouterWrapper_1_io_inChannels_3_credit_0_grant ),
       .io_inChannels_2_flit_x( CreditBuffer_2_io_out_2_flit_x ),
       .io_inChannels_2_flitValid( CreditBuffer_2_io_out_2_flitValid ),
       .io_inChannels_2_credit_1_grant( VCRouterWrapper_1_io_inChannels_2_credit_1_grant ),
       .io_inChannels_2_credit_0_grant( VCRouterWrapper_1_io_inChannels_2_credit_0_grant ),
       .io_inChannels_1_flit_x( CreditBuffer_io_out_1_flit_x ),
       .io_inChannels_1_flitValid( CreditBuffer_io_out_1_flitValid ),
       .io_inChannels_1_credit_1_grant( VCRouterWrapper_1_io_inChannels_1_credit_1_grant ),
       .io_inChannels_1_credit_0_grant( VCRouterWrapper_1_io_inChannels_1_credit_0_grant ),
       .io_inChannels_0_flit_x( io_inChannels_1_flit_x ),
       .io_inChannels_0_flitValid( io_inChannels_1_flitValid ),
       .io_inChannels_0_credit_1_grant( VCRouterWrapper_1_io_inChannels_0_credit_1_grant ),
       .io_inChannels_0_credit_0_grant( VCRouterWrapper_1_io_inChannels_0_credit_0_grant ),
       .io_outChannels_4_flit_x( VCRouterWrapper_1_io_outChannels_4_flit_x ),
       .io_outChannels_4_flitValid( VCRouterWrapper_1_io_outChannels_4_flitValid ),
       //.io_outChannels_4_credit_1_grant(  )
       //.io_outChannels_4_credit_0_grant(  )
       .io_outChannels_3_flit_x( VCRouterWrapper_1_io_outChannels_3_flit_x ),
       .io_outChannels_3_flitValid( VCRouterWrapper_1_io_outChannels_3_flitValid ),
       //.io_outChannels_3_credit_1_grant(  )
       //.io_outChannels_3_credit_0_grant(  )
       .io_outChannels_2_flit_x( VCRouterWrapper_1_io_outChannels_2_flit_x ),
       .io_outChannels_2_flitValid( VCRouterWrapper_1_io_outChannels_2_flitValid ),
       .io_outChannels_2_credit_1_grant( CreditBuffer_1_io_in_2_credit_1_grant ),
       .io_outChannels_2_credit_0_grant( CreditBuffer_1_io_in_2_credit_0_grant ),
       .io_outChannels_1_flit_x( VCRouterWrapper_1_io_outChannels_1_flit_x ),
       .io_outChannels_1_flitValid( VCRouterWrapper_1_io_outChannels_1_flitValid ),
       .io_outChannels_1_credit_1_grant( CreditBuffer_1_io_in_1_credit_1_grant ),
       .io_outChannels_1_credit_0_grant( CreditBuffer_1_io_in_1_credit_0_grant ),
       .io_outChannels_0_flit_x( VCRouterWrapper_1_io_outChannels_0_flit_x ),
       .io_outChannels_0_flitValid( VCRouterWrapper_1_io_outChannels_0_flitValid ),
       .io_outChannels_0_credit_1_grant( io_outChannels_1_credit_1_grant ),
       .io_outChannels_0_credit_0_grant( io_outChannels_1_credit_0_grant ),
       //.io_counters_1_counterVal(  )
       //.io_counters_1_counterIndex(  )
       //.io_counters_0_counterVal(  )
       //.io_counters_0_counterIndex(  )
       .io_bypass( io_bypass_1 )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign VCRouterWrapper_1.io_outChannels_4_credit_1_grant = {1{1'b0}};
    assign VCRouterWrapper_1.io_outChannels_4_credit_0_grant = {1{1'b0}};
    assign VCRouterWrapper_1.io_outChannels_3_credit_1_grant = {1{1'b0}};
    assign VCRouterWrapper_1.io_outChannels_3_credit_0_grant = {1{1'b0}};
// synthesis translate_on
`endif
  BusProbe_1 BusProbe_1(.clk(clk), .reset(reset),
       //.io_inFlit_4_x(  )
       //.io_inFlit_3_x(  )
       .io_inFlit_2_x( VCRouterWrapper_1_io_outChannels_2_flit_x ),
       .io_inFlit_1_x( VCRouterWrapper_1_io_outChannels_1_flit_x ),
       //.io_inFlit_0_x(  )
       //.io_inValid_4(  )
       //.io_inValid_3(  )
       .io_inValid_2( VCRouterWrapper_1_io_outChannels_2_flitValid ),
       .io_inValid_1( VCRouterWrapper_1_io_outChannels_1_flitValid ),
       //.io_inValid_0(  )
       .io_routerCord( 1'h0 ),
       //.io_startRecording(  )
       //.io_cyclesChannelBusy_4(  )
       //.io_cyclesChannelBusy_3(  )
       .io_cyclesChannelBusy_2( BusProbe_1_io_cyclesChannelBusy_2 ),
       .io_cyclesChannelBusy_1( BusProbe_1_io_cyclesChannelBusy_1 ),
       //.io_cyclesChannelBusy_0(  )
       .io_cyclesRouterBusy( BusProbe_1_io_cyclesRouterBusy )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign BusProbe_1.io_inValid_4 = {1{1'b0}};
    assign BusProbe_1.io_inValid_3 = {1{1'b0}};
    assign BusProbe_1.io_inValid_0 = {1{1'b0}};
// synthesis translate_on
`endif
  CreditBuffer CreditBuffer_1(.clk(clk), .reset(reset),
       //.io_in_4_flit_x(  )
       //.io_in_4_flitValid(  )
       //.io_in_4_credit_1_grant(  )
       //.io_in_4_credit_0_grant(  )
       //.io_in_3_flit_x(  )
       //.io_in_3_flitValid(  )
       //.io_in_3_credit_1_grant(  )
       //.io_in_3_credit_0_grant(  )
       .io_in_2_flit_x( VCRouterWrapper_1_io_outChannels_2_flit_x ),
       .io_in_2_flitValid( VCRouterWrapper_1_io_outChannels_2_flitValid ),
       .io_in_2_credit_1_grant( CreditBuffer_1_io_in_2_credit_1_grant ),
       .io_in_2_credit_0_grant( CreditBuffer_1_io_in_2_credit_0_grant ),
       .io_in_1_flit_x( VCRouterWrapper_1_io_outChannels_1_flit_x ),
       .io_in_1_flitValid( VCRouterWrapper_1_io_outChannels_1_flitValid ),
       .io_in_1_credit_1_grant( CreditBuffer_1_io_in_1_credit_1_grant ),
       .io_in_1_credit_0_grant( CreditBuffer_1_io_in_1_credit_0_grant ),
       //.io_in_0_flit_x(  )
       //.io_in_0_flitValid(  )
       //.io_in_0_credit_1_grant(  )
       //.io_in_0_credit_0_grant(  )
       //.io_out_4_flit_x(  )
       //.io_out_4_flitValid(  )
       //.io_out_4_credit_1_grant(  )
       //.io_out_4_credit_0_grant(  )
       //.io_out_3_flit_x(  )
       //.io_out_3_flitValid(  )
       //.io_out_3_credit_1_grant(  )
       //.io_out_3_credit_0_grant(  )
       .io_out_2_flit_x( CreditBuffer_1_io_out_2_flit_x ),
       .io_out_2_flitValid( CreditBuffer_1_io_out_2_flitValid ),
       .io_out_2_credit_1_grant( VCRouterWrapper_io_inChannels_2_credit_1_grant ),
       .io_out_2_credit_0_grant( VCRouterWrapper_io_inChannels_2_credit_0_grant ),
       .io_out_1_flit_x( CreditBuffer_1_io_out_1_flit_x ),
       .io_out_1_flitValid( CreditBuffer_1_io_out_1_flitValid ),
       .io_out_1_credit_1_grant( VCRouterWrapper_2_io_inChannels_1_credit_1_grant ),
       .io_out_1_credit_0_grant( VCRouterWrapper_2_io_inChannels_1_credit_0_grant )
       //.io_out_0_flit_x(  )
       //.io_out_0_flitValid(  )
       //.io_out_0_credit_1_grant(  )
       //.io_out_0_credit_0_grant(  )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign CreditBuffer_1.io_in_4_flit_x = {2{1'b0}};
    assign CreditBuffer_1.io_in_4_flitValid = {1{1'b0}};
    assign CreditBuffer_1.io_in_3_flit_x = {2{1'b0}};
    assign CreditBuffer_1.io_in_3_flitValid = {1{1'b0}};
    assign CreditBuffer_1.io_in_0_flit_x = {2{1'b0}};
    assign CreditBuffer_1.io_in_0_flitValid = {1{1'b0}};
    assign CreditBuffer_1.io_out_4_credit_1_grant = {1{1'b0}};
    assign CreditBuffer_1.io_out_4_credit_0_grant = {1{1'b0}};
    assign CreditBuffer_1.io_out_3_credit_1_grant = {1{1'b0}};
    assign CreditBuffer_1.io_out_3_credit_0_grant = {1{1'b0}};
    assign CreditBuffer_1.io_out_0_credit_1_grant = {1{1'b0}};
    assign CreditBuffer_1.io_out_0_credit_0_grant = {1{1'b0}};
// synthesis translate_on
`endif
  VCRouterWrapper_2 VCRouterWrapper_2(.clk(clk), .reset(reset),
       .io_inChannels_4_flit_x( OpenSoC_VCConstantEndpoint_7_io_outChannels_4_flit_x ),
       .io_inChannels_4_flitValid( OpenSoC_VCConstantEndpoint_7_io_outChannels_4_flitValid ),
       .io_inChannels_4_credit_1_grant( VCRouterWrapper_2_io_inChannels_4_credit_1_grant ),
       .io_inChannels_4_credit_0_grant( VCRouterWrapper_2_io_inChannels_4_credit_0_grant ),
       .io_inChannels_3_flit_x( OpenSoC_VCConstantEndpoint_6_io_outChannels_3_flit_x ),
       .io_inChannels_3_flitValid( OpenSoC_VCConstantEndpoint_6_io_outChannels_3_flitValid ),
       .io_inChannels_3_credit_1_grant( VCRouterWrapper_2_io_inChannels_3_credit_1_grant ),
       .io_inChannels_3_credit_0_grant( VCRouterWrapper_2_io_inChannels_3_credit_0_grant ),
       .io_inChannels_2_flit_x( OpenSoC_VCConstantEndpoint_5_io_outChannels_2_flit_x ),
       .io_inChannels_2_flitValid( OpenSoC_VCConstantEndpoint_5_io_outChannels_2_flitValid ),
       .io_inChannels_2_credit_1_grant( VCRouterWrapper_2_io_inChannels_2_credit_1_grant ),
       .io_inChannels_2_credit_0_grant( VCRouterWrapper_2_io_inChannels_2_credit_0_grant ),
       .io_inChannels_1_flit_x( CreditBuffer_1_io_out_1_flit_x ),
       .io_inChannels_1_flitValid( CreditBuffer_1_io_out_1_flitValid ),
       .io_inChannels_1_credit_1_grant( VCRouterWrapper_2_io_inChannels_1_credit_1_grant ),
       .io_inChannels_1_credit_0_grant( VCRouterWrapper_2_io_inChannels_1_credit_0_grant ),
       .io_inChannels_0_flit_x( io_inChannels_2_flit_x ),
       .io_inChannels_0_flitValid( io_inChannels_2_flitValid ),
       .io_inChannels_0_credit_1_grant( VCRouterWrapper_2_io_inChannels_0_credit_1_grant ),
       .io_inChannels_0_credit_0_grant( VCRouterWrapper_2_io_inChannels_0_credit_0_grant ),
       .io_outChannels_4_flit_x( VCRouterWrapper_2_io_outChannels_4_flit_x ),
       .io_outChannels_4_flitValid( VCRouterWrapper_2_io_outChannels_4_flitValid ),
       //.io_outChannels_4_credit_1_grant(  )
       //.io_outChannels_4_credit_0_grant(  )
       .io_outChannels_3_flit_x( VCRouterWrapper_2_io_outChannels_3_flit_x ),
       .io_outChannels_3_flitValid( VCRouterWrapper_2_io_outChannels_3_flitValid ),
       //.io_outChannels_3_credit_1_grant(  )
       //.io_outChannels_3_credit_0_grant(  )
       .io_outChannels_2_flit_x( VCRouterWrapper_2_io_outChannels_2_flit_x ),
       .io_outChannels_2_flitValid( VCRouterWrapper_2_io_outChannels_2_flitValid ),
       .io_outChannels_2_credit_1_grant( CreditBuffer_2_io_in_2_credit_1_grant ),
       .io_outChannels_2_credit_0_grant( CreditBuffer_2_io_in_2_credit_0_grant ),
       //.io_outChannels_1_flit_x(  )
       //.io_outChannels_1_flitValid(  )
       //.io_outChannels_1_credit_1_grant(  )
       //.io_outChannels_1_credit_0_grant(  )
       .io_outChannels_0_flit_x( VCRouterWrapper_2_io_outChannels_0_flit_x ),
       .io_outChannels_0_flitValid( VCRouterWrapper_2_io_outChannels_0_flitValid ),
       .io_outChannels_0_credit_1_grant( io_outChannels_2_credit_1_grant ),
       .io_outChannels_0_credit_0_grant( io_outChannels_2_credit_0_grant ),
       //.io_counters_1_counterVal(  )
       //.io_counters_1_counterIndex(  )
       //.io_counters_0_counterVal(  )
       //.io_counters_0_counterIndex(  )
       .io_bypass( io_bypass_2 )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign VCRouterWrapper_2.io_outChannels_4_credit_1_grant = {1{1'b0}};
    assign VCRouterWrapper_2.io_outChannels_4_credit_0_grant = {1{1'b0}};
    assign VCRouterWrapper_2.io_outChannels_3_credit_1_grant = {1{1'b0}};
    assign VCRouterWrapper_2.io_outChannels_3_credit_0_grant = {1{1'b0}};
    assign VCRouterWrapper_2.io_outChannels_1_credit_1_grant = {1{1'b0}};
    assign VCRouterWrapper_2.io_outChannels_1_credit_0_grant = {1{1'b0}};
// synthesis translate_on
`endif
  BusProbe_2 BusProbe_2(.clk(clk), .reset(reset),
       //.io_inFlit_4_x(  )
       //.io_inFlit_3_x(  )
       .io_inFlit_2_x( VCRouterWrapper_2_io_outChannels_2_flit_x ),
       //.io_inFlit_1_x(  )
       //.io_inFlit_0_x(  )
       //.io_inValid_4(  )
       //.io_inValid_3(  )
       .io_inValid_2( VCRouterWrapper_2_io_outChannels_2_flitValid ),
       //.io_inValid_1(  )
       //.io_inValid_0(  )
       .io_routerCord( 1'h0 ),
       //.io_startRecording(  )
       //.io_cyclesChannelBusy_4(  )
       //.io_cyclesChannelBusy_3(  )
       .io_cyclesChannelBusy_2( BusProbe_2_io_cyclesChannelBusy_2 ),
       //.io_cyclesChannelBusy_1(  )
       //.io_cyclesChannelBusy_0(  )
       .io_cyclesRouterBusy( BusProbe_2_io_cyclesRouterBusy )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign BusProbe_2.io_inValid_4 = {1{1'b0}};
    assign BusProbe_2.io_inValid_3 = {1{1'b0}};
    assign BusProbe_2.io_inValid_1 = {1{1'b0}};
    assign BusProbe_2.io_inValid_0 = {1{1'b0}};
// synthesis translate_on
`endif
  CreditBuffer CreditBuffer_2(.clk(clk), .reset(reset),
       //.io_in_4_flit_x(  )
       //.io_in_4_flitValid(  )
       //.io_in_4_credit_1_grant(  )
       //.io_in_4_credit_0_grant(  )
       //.io_in_3_flit_x(  )
       //.io_in_3_flitValid(  )
       //.io_in_3_credit_1_grant(  )
       //.io_in_3_credit_0_grant(  )
       .io_in_2_flit_x( VCRouterWrapper_2_io_outChannels_2_flit_x ),
       .io_in_2_flitValid( VCRouterWrapper_2_io_outChannels_2_flitValid ),
       .io_in_2_credit_1_grant( CreditBuffer_2_io_in_2_credit_1_grant ),
       .io_in_2_credit_0_grant( CreditBuffer_2_io_in_2_credit_0_grant ),
       //.io_in_1_flit_x(  )
       //.io_in_1_flitValid(  )
       //.io_in_1_credit_1_grant(  )
       //.io_in_1_credit_0_grant(  )
       //.io_in_0_flit_x(  )
       //.io_in_0_flitValid(  )
       //.io_in_0_credit_1_grant(  )
       //.io_in_0_credit_0_grant(  )
       //.io_out_4_flit_x(  )
       //.io_out_4_flitValid(  )
       //.io_out_4_credit_1_grant(  )
       //.io_out_4_credit_0_grant(  )
       //.io_out_3_flit_x(  )
       //.io_out_3_flitValid(  )
       //.io_out_3_credit_1_grant(  )
       //.io_out_3_credit_0_grant(  )
       .io_out_2_flit_x( CreditBuffer_2_io_out_2_flit_x ),
       .io_out_2_flitValid( CreditBuffer_2_io_out_2_flitValid ),
       .io_out_2_credit_1_grant( VCRouterWrapper_1_io_inChannels_2_credit_1_grant ),
       .io_out_2_credit_0_grant( VCRouterWrapper_1_io_inChannels_2_credit_0_grant )
       //.io_out_1_flit_x(  )
       //.io_out_1_flitValid(  )
       //.io_out_1_credit_1_grant(  )
       //.io_out_1_credit_0_grant(  )
       //.io_out_0_flit_x(  )
       //.io_out_0_flitValid(  )
       //.io_out_0_credit_1_grant(  )
       //.io_out_0_credit_0_grant(  )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign CreditBuffer_2.io_in_4_flit_x = {2{1'b0}};
    assign CreditBuffer_2.io_in_4_flitValid = {1{1'b0}};
    assign CreditBuffer_2.io_in_3_flit_x = {2{1'b0}};
    assign CreditBuffer_2.io_in_3_flitValid = {1{1'b0}};
    assign CreditBuffer_2.io_in_1_flit_x = {2{1'b0}};
    assign CreditBuffer_2.io_in_1_flitValid = {1{1'b0}};
    assign CreditBuffer_2.io_in_0_flit_x = {2{1'b0}};
    assign CreditBuffer_2.io_in_0_flitValid = {1{1'b0}};
    assign CreditBuffer_2.io_out_4_credit_1_grant = {1{1'b0}};
    assign CreditBuffer_2.io_out_4_credit_0_grant = {1{1'b0}};
    assign CreditBuffer_2.io_out_3_credit_1_grant = {1{1'b0}};
    assign CreditBuffer_2.io_out_3_credit_0_grant = {1{1'b0}};
    assign CreditBuffer_2.io_out_1_credit_1_grant = {1{1'b0}};
    assign CreditBuffer_2.io_out_1_credit_0_grant = {1{1'b0}};
    assign CreditBuffer_2.io_out_0_credit_1_grant = {1{1'b0}};
    assign CreditBuffer_2.io_out_0_credit_0_grant = {1{1'b0}};
// synthesis translate_on
`endif
  OpenSoC_VCConstantEndpoint_0 OpenSoC_VCConstantEndpoint(
       //.io_inChannels_4_flit_x(  )
       //.io_inChannels_4_flitValid(  )
       //.io_inChannels_4_credit_1_grant(  )
       //.io_inChannels_4_credit_0_grant(  )
       //.io_inChannels_3_flit_x(  )
       //.io_inChannels_3_flitValid(  )
       //.io_inChannels_3_credit_1_grant(  )
       //.io_inChannels_3_credit_0_grant(  )
       //.io_inChannels_2_flit_x(  )
       //.io_inChannels_2_flitValid(  )
       //.io_inChannels_2_credit_1_grant(  )
       //.io_inChannels_2_credit_0_grant(  )
       .io_inChannels_1_flit_x( VCRouterWrapper_io_outChannels_1_flit_x ),
       .io_inChannels_1_flitValid( VCRouterWrapper_io_outChannels_1_flitValid ),
       //.io_inChannels_1_credit_1_grant(  )
       //.io_inChannels_1_credit_0_grant(  )
       //.io_inChannels_0_flit_x(  )
       //.io_inChannels_0_flitValid(  )
       //.io_inChannels_0_credit_1_grant(  )
       //.io_inChannels_0_credit_0_grant(  )
       //.io_outChannels_4_flit_x(  )
       //.io_outChannels_4_flitValid(  )
       //.io_outChannels_4_credit_1_grant(  )
       //.io_outChannels_4_credit_0_grant(  )
       //.io_outChannels_3_flit_x(  )
       //.io_outChannels_3_flitValid(  )
       //.io_outChannels_3_credit_1_grant(  )
       //.io_outChannels_3_credit_0_grant(  )
       //.io_outChannels_2_flit_x(  )
       //.io_outChannels_2_flitValid(  )
       //.io_outChannels_2_credit_1_grant(  )
       //.io_outChannels_2_credit_0_grant(  )
       .io_outChannels_1_flit_x( OpenSoC_VCConstantEndpoint_io_outChannels_1_flit_x ),
       .io_outChannels_1_flitValid( OpenSoC_VCConstantEndpoint_io_outChannels_1_flitValid ),
       .io_outChannels_1_credit_1_grant( VCRouterWrapper_io_inChannels_1_credit_1_grant ),
       .io_outChannels_1_credit_0_grant( VCRouterWrapper_io_inChannels_1_credit_0_grant )
       //.io_outChannels_0_flit_x(  )
       //.io_outChannels_0_flitValid(  )
       //.io_outChannels_0_credit_1_grant(  )
       //.io_outChannels_0_credit_0_grant(  )
       //.io_counters_1_counterVal(  )
       //.io_counters_1_counterIndex(  )
       //.io_counters_0_counterVal(  )
       //.io_counters_0_counterIndex(  )
       //.io_bypass(  )
  );
  OpenSoC_VCConstantEndpoint_1 OpenSoC_VCConstantEndpoint_1(
       //.io_inChannels_4_flit_x(  )
       //.io_inChannels_4_flitValid(  )
       //.io_inChannels_4_credit_1_grant(  )
       //.io_inChannels_4_credit_0_grant(  )
       .io_inChannels_3_flit_x( VCRouterWrapper_io_outChannels_3_flit_x ),
       .io_inChannels_3_flitValid( VCRouterWrapper_io_outChannels_3_flitValid ),
       //.io_inChannels_3_credit_1_grant(  )
       //.io_inChannels_3_credit_0_grant(  )
       //.io_inChannels_2_flit_x(  )
       //.io_inChannels_2_flitValid(  )
       //.io_inChannels_2_credit_1_grant(  )
       //.io_inChannels_2_credit_0_grant(  )
       //.io_inChannels_1_flit_x(  )
       //.io_inChannels_1_flitValid(  )
       //.io_inChannels_1_credit_1_grant(  )
       //.io_inChannels_1_credit_0_grant(  )
       //.io_inChannels_0_flit_x(  )
       //.io_inChannels_0_flitValid(  )
       //.io_inChannels_0_credit_1_grant(  )
       //.io_inChannels_0_credit_0_grant(  )
       //.io_outChannels_4_flit_x(  )
       //.io_outChannels_4_flitValid(  )
       //.io_outChannels_4_credit_1_grant(  )
       //.io_outChannels_4_credit_0_grant(  )
       .io_outChannels_3_flit_x( OpenSoC_VCConstantEndpoint_1_io_outChannels_3_flit_x ),
       .io_outChannels_3_flitValid( OpenSoC_VCConstantEndpoint_1_io_outChannels_3_flitValid ),
       .io_outChannels_3_credit_1_grant( VCRouterWrapper_io_inChannels_3_credit_1_grant ),
       .io_outChannels_3_credit_0_grant( VCRouterWrapper_io_inChannels_3_credit_0_grant )
       //.io_outChannels_2_flit_x(  )
       //.io_outChannels_2_flitValid(  )
       //.io_outChannels_2_credit_1_grant(  )
       //.io_outChannels_2_credit_0_grant(  )
       //.io_outChannels_1_flit_x(  )
       //.io_outChannels_1_flitValid(  )
       //.io_outChannels_1_credit_1_grant(  )
       //.io_outChannels_1_credit_0_grant(  )
       //.io_outChannels_0_flit_x(  )
       //.io_outChannels_0_flitValid(  )
       //.io_outChannels_0_credit_1_grant(  )
       //.io_outChannels_0_credit_0_grant(  )
       //.io_counters_1_counterVal(  )
       //.io_counters_1_counterIndex(  )
       //.io_counters_0_counterVal(  )
       //.io_counters_0_counterIndex(  )
       //.io_bypass(  )
  );
  OpenSoC_VCConstantEndpoint_2 OpenSoC_VCConstantEndpoint_2(
       .io_inChannels_4_flit_x( VCRouterWrapper_io_outChannels_4_flit_x ),
       .io_inChannels_4_flitValid( VCRouterWrapper_io_outChannels_4_flitValid ),
       //.io_inChannels_4_credit_1_grant(  )
       //.io_inChannels_4_credit_0_grant(  )
       //.io_inChannels_3_flit_x(  )
       //.io_inChannels_3_flitValid(  )
       //.io_inChannels_3_credit_1_grant(  )
       //.io_inChannels_3_credit_0_grant(  )
       //.io_inChannels_2_flit_x(  )
       //.io_inChannels_2_flitValid(  )
       //.io_inChannels_2_credit_1_grant(  )
       //.io_inChannels_2_credit_0_grant(  )
       //.io_inChannels_1_flit_x(  )
       //.io_inChannels_1_flitValid(  )
       //.io_inChannels_1_credit_1_grant(  )
       //.io_inChannels_1_credit_0_grant(  )
       //.io_inChannels_0_flit_x(  )
       //.io_inChannels_0_flitValid(  )
       //.io_inChannels_0_credit_1_grant(  )
       //.io_inChannels_0_credit_0_grant(  )
       .io_outChannels_4_flit_x( OpenSoC_VCConstantEndpoint_2_io_outChannels_4_flit_x ),
       .io_outChannels_4_flitValid( OpenSoC_VCConstantEndpoint_2_io_outChannels_4_flitValid ),
       .io_outChannels_4_credit_1_grant( VCRouterWrapper_io_inChannels_4_credit_1_grant ),
       .io_outChannels_4_credit_0_grant( VCRouterWrapper_io_inChannels_4_credit_0_grant )
       //.io_outChannels_3_flit_x(  )
       //.io_outChannels_3_flitValid(  )
       //.io_outChannels_3_credit_1_grant(  )
       //.io_outChannels_3_credit_0_grant(  )
       //.io_outChannels_2_flit_x(  )
       //.io_outChannels_2_flitValid(  )
       //.io_outChannels_2_credit_1_grant(  )
       //.io_outChannels_2_credit_0_grant(  )
       //.io_outChannels_1_flit_x(  )
       //.io_outChannels_1_flitValid(  )
       //.io_outChannels_1_credit_1_grant(  )
       //.io_outChannels_1_credit_0_grant(  )
       //.io_outChannels_0_flit_x(  )
       //.io_outChannels_0_flitValid(  )
       //.io_outChannels_0_credit_1_grant(  )
       //.io_outChannels_0_credit_0_grant(  )
       //.io_counters_1_counterVal(  )
       //.io_counters_1_counterIndex(  )
       //.io_counters_0_counterVal(  )
       //.io_counters_0_counterIndex(  )
       //.io_bypass(  )
  );
  OpenSoC_VCConstantEndpoint_1 OpenSoC_VCConstantEndpoint_3(
       //.io_inChannels_4_flit_x(  )
       //.io_inChannels_4_flitValid(  )
       //.io_inChannels_4_credit_1_grant(  )
       //.io_inChannels_4_credit_0_grant(  )
       .io_inChannels_3_flit_x( VCRouterWrapper_1_io_outChannels_3_flit_x ),
       .io_inChannels_3_flitValid( VCRouterWrapper_1_io_outChannels_3_flitValid ),
       //.io_inChannels_3_credit_1_grant(  )
       //.io_inChannels_3_credit_0_grant(  )
       //.io_inChannels_2_flit_x(  )
       //.io_inChannels_2_flitValid(  )
       //.io_inChannels_2_credit_1_grant(  )
       //.io_inChannels_2_credit_0_grant(  )
       //.io_inChannels_1_flit_x(  )
       //.io_inChannels_1_flitValid(  )
       //.io_inChannels_1_credit_1_grant(  )
       //.io_inChannels_1_credit_0_grant(  )
       //.io_inChannels_0_flit_x(  )
       //.io_inChannels_0_flitValid(  )
       //.io_inChannels_0_credit_1_grant(  )
       //.io_inChannels_0_credit_0_grant(  )
       //.io_outChannels_4_flit_x(  )
       //.io_outChannels_4_flitValid(  )
       //.io_outChannels_4_credit_1_grant(  )
       //.io_outChannels_4_credit_0_grant(  )
       .io_outChannels_3_flit_x( OpenSoC_VCConstantEndpoint_3_io_outChannels_3_flit_x ),
       .io_outChannels_3_flitValid( OpenSoC_VCConstantEndpoint_3_io_outChannels_3_flitValid ),
       .io_outChannels_3_credit_1_grant( VCRouterWrapper_1_io_inChannels_3_credit_1_grant ),
       .io_outChannels_3_credit_0_grant( VCRouterWrapper_1_io_inChannels_3_credit_0_grant )
       //.io_outChannels_2_flit_x(  )
       //.io_outChannels_2_flitValid(  )
       //.io_outChannels_2_credit_1_grant(  )
       //.io_outChannels_2_credit_0_grant(  )
       //.io_outChannels_1_flit_x(  )
       //.io_outChannels_1_flitValid(  )
       //.io_outChannels_1_credit_1_grant(  )
       //.io_outChannels_1_credit_0_grant(  )
       //.io_outChannels_0_flit_x(  )
       //.io_outChannels_0_flitValid(  )
       //.io_outChannels_0_credit_1_grant(  )
       //.io_outChannels_0_credit_0_grant(  )
       //.io_counters_1_counterVal(  )
       //.io_counters_1_counterIndex(  )
       //.io_counters_0_counterVal(  )
       //.io_counters_0_counterIndex(  )
       //.io_bypass(  )
  );
  OpenSoC_VCConstantEndpoint_2 OpenSoC_VCConstantEndpoint_4(
       .io_inChannels_4_flit_x( VCRouterWrapper_1_io_outChannels_4_flit_x ),
       .io_inChannels_4_flitValid( VCRouterWrapper_1_io_outChannels_4_flitValid ),
       //.io_inChannels_4_credit_1_grant(  )
       //.io_inChannels_4_credit_0_grant(  )
       //.io_inChannels_3_flit_x(  )
       //.io_inChannels_3_flitValid(  )
       //.io_inChannels_3_credit_1_grant(  )
       //.io_inChannels_3_credit_0_grant(  )
       //.io_inChannels_2_flit_x(  )
       //.io_inChannels_2_flitValid(  )
       //.io_inChannels_2_credit_1_grant(  )
       //.io_inChannels_2_credit_0_grant(  )
       //.io_inChannels_1_flit_x(  )
       //.io_inChannels_1_flitValid(  )
       //.io_inChannels_1_credit_1_grant(  )
       //.io_inChannels_1_credit_0_grant(  )
       //.io_inChannels_0_flit_x(  )
       //.io_inChannels_0_flitValid(  )
       //.io_inChannels_0_credit_1_grant(  )
       //.io_inChannels_0_credit_0_grant(  )
       .io_outChannels_4_flit_x( OpenSoC_VCConstantEndpoint_4_io_outChannels_4_flit_x ),
       .io_outChannels_4_flitValid( OpenSoC_VCConstantEndpoint_4_io_outChannels_4_flitValid ),
       .io_outChannels_4_credit_1_grant( VCRouterWrapper_1_io_inChannels_4_credit_1_grant ),
       .io_outChannels_4_credit_0_grant( VCRouterWrapper_1_io_inChannels_4_credit_0_grant )
       //.io_outChannels_3_flit_x(  )
       //.io_outChannels_3_flitValid(  )
       //.io_outChannels_3_credit_1_grant(  )
       //.io_outChannels_3_credit_0_grant(  )
       //.io_outChannels_2_flit_x(  )
       //.io_outChannels_2_flitValid(  )
       //.io_outChannels_2_credit_1_grant(  )
       //.io_outChannels_2_credit_0_grant(  )
       //.io_outChannels_1_flit_x(  )
       //.io_outChannels_1_flitValid(  )
       //.io_outChannels_1_credit_1_grant(  )
       //.io_outChannels_1_credit_0_grant(  )
       //.io_outChannels_0_flit_x(  )
       //.io_outChannels_0_flitValid(  )
       //.io_outChannels_0_credit_1_grant(  )
       //.io_outChannels_0_credit_0_grant(  )
       //.io_counters_1_counterVal(  )
       //.io_counters_1_counterIndex(  )
       //.io_counters_0_counterVal(  )
       //.io_counters_0_counterIndex(  )
       //.io_bypass(  )
  );
  OpenSoC_VCConstantEndpoint_3 OpenSoC_VCConstantEndpoint_5(
       //.io_inChannels_4_flit_x(  )
       //.io_inChannels_4_flitValid(  )
       //.io_inChannels_4_credit_1_grant(  )
       //.io_inChannels_4_credit_0_grant(  )
       //.io_inChannels_3_flit_x(  )
       //.io_inChannels_3_flitValid(  )
       //.io_inChannels_3_credit_1_grant(  )
       //.io_inChannels_3_credit_0_grant(  )
       .io_inChannels_2_flit_x( VCRouterWrapper_2_io_outChannels_2_flit_x ),
       .io_inChannels_2_flitValid( VCRouterWrapper_2_io_outChannels_2_flitValid ),
       //.io_inChannels_2_credit_1_grant(  )
       //.io_inChannels_2_credit_0_grant(  )
       //.io_inChannels_1_flit_x(  )
       //.io_inChannels_1_flitValid(  )
       //.io_inChannels_1_credit_1_grant(  )
       //.io_inChannels_1_credit_0_grant(  )
       //.io_inChannels_0_flit_x(  )
       //.io_inChannels_0_flitValid(  )
       //.io_inChannels_0_credit_1_grant(  )
       //.io_inChannels_0_credit_0_grant(  )
       //.io_outChannels_4_flit_x(  )
       //.io_outChannels_4_flitValid(  )
       //.io_outChannels_4_credit_1_grant(  )
       //.io_outChannels_4_credit_0_grant(  )
       //.io_outChannels_3_flit_x(  )
       //.io_outChannels_3_flitValid(  )
       //.io_outChannels_3_credit_1_grant(  )
       //.io_outChannels_3_credit_0_grant(  )
       .io_outChannels_2_flit_x( OpenSoC_VCConstantEndpoint_5_io_outChannels_2_flit_x ),
       .io_outChannels_2_flitValid( OpenSoC_VCConstantEndpoint_5_io_outChannels_2_flitValid ),
       .io_outChannels_2_credit_1_grant( VCRouterWrapper_2_io_inChannels_2_credit_1_grant ),
       .io_outChannels_2_credit_0_grant( VCRouterWrapper_2_io_inChannels_2_credit_0_grant )
       //.io_outChannels_1_flit_x(  )
       //.io_outChannels_1_flitValid(  )
       //.io_outChannels_1_credit_1_grant(  )
       //.io_outChannels_1_credit_0_grant(  )
       //.io_outChannels_0_flit_x(  )
       //.io_outChannels_0_flitValid(  )
       //.io_outChannels_0_credit_1_grant(  )
       //.io_outChannels_0_credit_0_grant(  )
       //.io_counters_1_counterVal(  )
       //.io_counters_1_counterIndex(  )
       //.io_counters_0_counterVal(  )
       //.io_counters_0_counterIndex(  )
       //.io_bypass(  )
  );
  OpenSoC_VCConstantEndpoint_1 OpenSoC_VCConstantEndpoint_6(
       //.io_inChannels_4_flit_x(  )
       //.io_inChannels_4_flitValid(  )
       //.io_inChannels_4_credit_1_grant(  )
       //.io_inChannels_4_credit_0_grant(  )
       .io_inChannels_3_flit_x( VCRouterWrapper_2_io_outChannels_3_flit_x ),
       .io_inChannels_3_flitValid( VCRouterWrapper_2_io_outChannels_3_flitValid ),
       //.io_inChannels_3_credit_1_grant(  )
       //.io_inChannels_3_credit_0_grant(  )
       //.io_inChannels_2_flit_x(  )
       //.io_inChannels_2_flitValid(  )
       //.io_inChannels_2_credit_1_grant(  )
       //.io_inChannels_2_credit_0_grant(  )
       //.io_inChannels_1_flit_x(  )
       //.io_inChannels_1_flitValid(  )
       //.io_inChannels_1_credit_1_grant(  )
       //.io_inChannels_1_credit_0_grant(  )
       //.io_inChannels_0_flit_x(  )
       //.io_inChannels_0_flitValid(  )
       //.io_inChannels_0_credit_1_grant(  )
       //.io_inChannels_0_credit_0_grant(  )
       //.io_outChannels_4_flit_x(  )
       //.io_outChannels_4_flitValid(  )
       //.io_outChannels_4_credit_1_grant(  )
       //.io_outChannels_4_credit_0_grant(  )
       .io_outChannels_3_flit_x( OpenSoC_VCConstantEndpoint_6_io_outChannels_3_flit_x ),
       .io_outChannels_3_flitValid( OpenSoC_VCConstantEndpoint_6_io_outChannels_3_flitValid ),
       .io_outChannels_3_credit_1_grant( VCRouterWrapper_2_io_inChannels_3_credit_1_grant ),
       .io_outChannels_3_credit_0_grant( VCRouterWrapper_2_io_inChannels_3_credit_0_grant )
       //.io_outChannels_2_flit_x(  )
       //.io_outChannels_2_flitValid(  )
       //.io_outChannels_2_credit_1_grant(  )
       //.io_outChannels_2_credit_0_grant(  )
       //.io_outChannels_1_flit_x(  )
       //.io_outChannels_1_flitValid(  )
       //.io_outChannels_1_credit_1_grant(  )
       //.io_outChannels_1_credit_0_grant(  )
       //.io_outChannels_0_flit_x(  )
       //.io_outChannels_0_flitValid(  )
       //.io_outChannels_0_credit_1_grant(  )
       //.io_outChannels_0_credit_0_grant(  )
       //.io_counters_1_counterVal(  )
       //.io_counters_1_counterIndex(  )
       //.io_counters_0_counterVal(  )
       //.io_counters_0_counterIndex(  )
       //.io_bypass(  )
  );
  OpenSoC_VCConstantEndpoint_2 OpenSoC_VCConstantEndpoint_7(
       .io_inChannels_4_flit_x( VCRouterWrapper_2_io_outChannels_4_flit_x ),
       .io_inChannels_4_flitValid( VCRouterWrapper_2_io_outChannels_4_flitValid ),
       //.io_inChannels_4_credit_1_grant(  )
       //.io_inChannels_4_credit_0_grant(  )
       //.io_inChannels_3_flit_x(  )
       //.io_inChannels_3_flitValid(  )
       //.io_inChannels_3_credit_1_grant(  )
       //.io_inChannels_3_credit_0_grant(  )
       //.io_inChannels_2_flit_x(  )
       //.io_inChannels_2_flitValid(  )
       //.io_inChannels_2_credit_1_grant(  )
       //.io_inChannels_2_credit_0_grant(  )
       //.io_inChannels_1_flit_x(  )
       //.io_inChannels_1_flitValid(  )
       //.io_inChannels_1_credit_1_grant(  )
       //.io_inChannels_1_credit_0_grant(  )
       //.io_inChannels_0_flit_x(  )
       //.io_inChannels_0_flitValid(  )
       //.io_inChannels_0_credit_1_grant(  )
       //.io_inChannels_0_credit_0_grant(  )
       .io_outChannels_4_flit_x( OpenSoC_VCConstantEndpoint_7_io_outChannels_4_flit_x ),
       .io_outChannels_4_flitValid( OpenSoC_VCConstantEndpoint_7_io_outChannels_4_flitValid ),
       .io_outChannels_4_credit_1_grant( VCRouterWrapper_2_io_inChannels_4_credit_1_grant ),
       .io_outChannels_4_credit_0_grant( VCRouterWrapper_2_io_inChannels_4_credit_0_grant )
       //.io_outChannels_3_flit_x(  )
       //.io_outChannels_3_flitValid(  )
       //.io_outChannels_3_credit_1_grant(  )
       //.io_outChannels_3_credit_0_grant(  )
       //.io_outChannels_2_flit_x(  )
       //.io_outChannels_2_flitValid(  )
       //.io_outChannels_2_credit_1_grant(  )
       //.io_outChannels_2_credit_0_grant(  )
       //.io_outChannels_1_flit_x(  )
       //.io_outChannels_1_flitValid(  )
       //.io_outChannels_1_credit_1_grant(  )
       //.io_outChannels_1_credit_0_grant(  )
       //.io_outChannels_0_flit_x(  )
       //.io_outChannels_0_flitValid(  )
       //.io_outChannels_0_credit_1_grant(  )
       //.io_outChannels_0_credit_0_grant(  )
       //.io_counters_1_counterVal(  )
       //.io_counters_1_counterIndex(  )
       //.io_counters_0_counterVal(  )
       //.io_counters_0_counterIndex(  )
       //.io_bypass(  )
  );
endmodule

module RRArbiter_0(input clk, input reset,
    input  io_requests_1_releaseLock,
    output io_requests_1_grant,
    input  io_requests_1_request,
    //input [2:0] io_requests_1_priorityLevel
    input  io_requests_0_releaseLock,
    output io_requests_0_grant,
    input  io_requests_0_request,
    //input [2:0] io_requests_0_priorityLevel
    input  io_resource_ready,
    output io_resource_valid,
    output io_chosen
);

  wire T53;
  wire[1:0] winner;
  wire[1:0] T1;
  reg [1:0] nextGrant;
  wire[1:0] T54;
  wire[1:0] T2;
  wire[1:0] T3;
  wire T4;
  wire[1:0] T5;
  wire[1:0] requestsBits;
  wire T6;
  wire T7;
  wire[1:0] T8;
  wire[1:0] T9;
  wire[2:0] passSelectL0;
  wire[2:0] T10;
  wire[2:0] T11;
  wire[2:0] T12;
  wire[1:0] T13;
  wire T14;
  wire T15;
  wire T16;
  wire[2:0] T17;
  wire[1:0] T18;
  wire T19;
  wire[1:0] passSelectL1;
  wire[1:0] T20;
  wire[1:0] T21;
  wire[1:0] T55;
  wire T22;
  wire[1:0] T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire lockRelease;
  wire T28;
  wire T29;
  wire nextGrantUInt;
  wire T56;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  wire T52;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    nextGrant = {1{1'b0}};
  end
// synthesis translate_on
`endif

  assign io_chosen = T53;
  assign T53 = winner[1'h1:1'h1];
  assign winner = T1;
  assign T1 = T25 ? T5 : nextGrant;
  assign T54 = reset ? 2'h2 : T2;
  assign T2 = T25 ? T3 : nextGrant;
  assign T3 = T4 ? winner : nextGrant;
  assign T4 = winner != 2'h0;
  assign T5 = T8 & requestsBits;
  assign requestsBits = {T7, T6};
  assign T6 = io_requests_0_request;
  assign T7 = io_requests_1_request;
  assign T8 = T24 ? passSelectL1 : T9;
  assign T9 = passSelectL0[1'h1:1'h0];
  assign passSelectL0 = T10;
  assign T10 = T25 ? T11 : 3'h0;
  assign T11 = T17 + T12;
  assign T12 = {T16, T13};
  assign T13 = {T15, T14};
  assign T14 = nextGrant[1'h1:1'h1];
  assign T15 = nextGrant[1'h0:1'h0];
  assign T16 = 1'h0;
  assign T17 = {T19, T18};
  assign T18 = ~ requestsBits;
  assign T19 = 1'h0;
  assign passSelectL1 = T20;
  assign T20 = T25 ? T21 : 2'h0;
  assign T21 = T23 + T55;
  assign T55 = {1'h0, T22};
  assign T22 = 1'h1;
  assign T23 = ~ requestsBits;
  assign T24 = passSelectL0[2'h2:2'h2];
  assign T25 = T26 ^ 1'h1;
  assign T26 = T31 & T27;
  assign T27 = ~ lockRelease;
  assign lockRelease = T28;
  assign T28 = T29 ? io_requests_1_releaseLock : io_requests_0_releaseLock;
  assign T29 = nextGrantUInt;
  assign nextGrantUInt = T56;
  assign T56 = nextGrant[1'h1:1'h1];
  assign T31 = T38 & T32;
  assign T32 = T37 & T33;
  assign T33 = T34 - 1'h1;
  assign T34 = 1'h1 << T35;
  assign T35 = T36 + 1'h1;
  assign T36 = nextGrantUInt - nextGrantUInt;
  assign T37 = requestsBits >> nextGrantUInt;
  assign T38 = T43 & T39;
  assign T39 = T40 - 1'h1;
  assign T40 = 1'h1 << T41;
  assign T41 = T42 + 1'h1;
  assign T42 = nextGrantUInt - nextGrantUInt;
  assign T43 = nextGrant >> nextGrantUInt;
  assign io_resource_valid = T44;
  assign T44 = T45 & io_resource_ready;
  assign T45 = T46 ? io_requests_1_grant : io_requests_0_grant;
  assign T46 = io_chosen;
  assign io_requests_0_grant = T47;
  assign T47 = T48 & io_resource_ready;
  assign T48 = T49;
  assign T49 = winner[1'h0:1'h0];
  assign io_requests_1_grant = T50;
  assign T50 = T51 & io_resource_ready;
  assign T51 = T52;
  assign T52 = winner[1'h1:1'h1];

  always @(posedge clk) begin
    if(reset) begin
      nextGrant <= 2'h2;
    end else if(T25) begin
      nextGrant <= T3;
    end
  end
endmodule

module InjectionQStateMgmt(input clk, input reset,
    input  io_inputBufferValid,
    input  io_creditsAvailable,
    input  io_inputIsTail,
    input  io_vcAllocGranted,
    output[1:0] io_currentState
);

  reg [1:0] curState;
  wire[1:0] T38;
  wire[1:0] T0;
  wire[1:0] T1;
  wire[1:0] T2;
  wire[1:0] T3;
  wire[1:0] T4;
  wire[1:0] T5;
  wire[1:0] T6;
  wire[1:0] T7;
  wire[1:0] T8;
  wire T9;
  wire T10;
  wire T11;
  wire T12;
  wire T13;
  wire T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    curState = {1{1'b0}};
  end
// synthesis translate_on
`endif

  assign io_currentState = curState;
  assign T38 = reset ? 2'h0 : T0;
  assign T0 = T36 ? 2'h3 : T1;
  assign T1 = T31 ? 2'h2 : T2;
  assign T2 = T29 ? 2'h2 : T3;
  assign T3 = T26 ? 2'h0 : T4;
  assign T4 = T20 ? 2'h3 : T5;
  assign T5 = T18 ? 2'h1 : T6;
  assign T6 = T14 ? 2'h2 : T7;
  assign T7 = T12 ? 2'h0 : T8;
  assign T8 = T9 ? 2'h1 : curState;
  assign T9 = T11 & T10;
  assign T10 = io_inputBufferValid & io_vcAllocGranted;
  assign T11 = curState == 2'h0;
  assign T12 = T11 & T13;
  assign T13 = T10 ^ 1'h1;
  assign T14 = T15 & io_creditsAvailable;
  assign T15 = T17 & T16;
  assign T16 = curState == 2'h1;
  assign T17 = T11 ^ 1'h1;
  assign T18 = T15 & T19;
  assign T19 = io_creditsAvailable ^ 1'h1;
  assign T20 = T22 & T21;
  assign T21 = io_creditsAvailable ^ 1'h1;
  assign T22 = T24 & T23;
  assign T23 = curState == 2'h2;
  assign T24 = T25 ^ 1'h1;
  assign T25 = T11 | T16;
  assign T26 = T27 & io_inputIsTail;
  assign T27 = T22 & T28;
  assign T28 = T21 ^ 1'h1;
  assign T29 = T27 & T30;
  assign T30 = io_inputIsTail ^ 1'h1;
  assign T31 = T32 & io_creditsAvailable;
  assign T32 = T34 & T33;
  assign T33 = curState == 2'h3;
  assign T34 = T35 ^ 1'h1;
  assign T35 = T25 | T23;
  assign T36 = T32 & T37;
  assign T37 = io_creditsAvailable ^ 1'h1;

  always @(posedge clk) begin
    if(reset) begin
      curState <= 2'h0;
    end else if(T36) begin
      curState <= 2'h3;
    end else if(T31) begin
      curState <= 2'h2;
    end else if(T29) begin
      curState <= 2'h2;
    end else if(T26) begin
      curState <= 2'h0;
    end else if(T20) begin
      curState <= 2'h3;
    end else if(T18) begin
      curState <= 2'h1;
    end else if(T14) begin
      curState <= 2'h2;
    end else if(T12) begin
      curState <= 2'h0;
    end else if(T9) begin
      curState <= 2'h1;
    end
  end
endmodule

module InjectionChannelQ(input clk, input reset,
    input [54:0] io_in_flit_x,
    input  io_in_flitValid,
    output io_in_credit_grant,
    output[54:0] io_out_flit_x,
    output io_out_flitValid,
    input  io_out_credit_1_grant,
    input  io_out_credit_0_grant
);

  wire T0;
  wire T1;
  wire T2;
  wire T3;
  wire T4;
  wire T5;
  wire T6;
  wire[4:0] T7;
  wire T8;
  wire T9;
  wire T10;
  wire T11;
  wire[53:0] T12;
  wire T13;
  wire[30:0] T14;
  wire T15;
  wire T16;
  wire T17;
  wire T18;
  wire T19;
  wire T20;
  wire T21;
  wire T22;
  wire T23;
  wire T24;
  wire T25;
  wire T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  wire T32;
  wire T33;
  wire T34;
  wire T35;
  wire T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire creditGen_io_outCredit_grant;
  wire CreditCon_io_outCredit;
  wire CreditCon_io_almostOut;
  wire CreditCon_1_io_outCredit;
  wire CreditCon_1_io_almostOut;
  wire vcArbiter_io_requests_1_grant;
  wire vcArbiter_io_requests_0_grant;
  wire vcArbiter_io_resource_valid;
  wire vcArbiter_io_chosen;
  wire[1:0] injQStateMachine_io_currentState;
  wire queue_io_deq_valid;
  wire[54:0] queue_io_deq_bits_x;
  wire[4:0] queue_io_count;
  wire[54:0] replaceVC_io_newFlit_x;


  assign T0 = T2 & T1;
  assign T1 = injQStateMachine_io_currentState == 2'h2;
  assign T2 = T3 & vcArbiter_io_resource_valid;
  assign T3 = T4 ? CreditCon_1_io_outCredit : CreditCon_io_outCredit;
  assign T4 = vcArbiter_io_chosen;
  assign T5 = T6 & io_in_flitValid;
  assign T6 = 5'h1 < T7;
  assign T7 = 5'h10 - queue_io_count;
  assign T8 = T9 & queue_io_deq_valid;
  assign T9 = T10;
  assign T10 = T15 ? T13 : T11;
  assign T11 = T12[6'h25:6'h25];
  assign T12 = queue_io_deq_bits_x[6'h36:1'h1];
  assign T13 = T14[4'he:4'he];
  assign T14 = queue_io_deq_bits_x[5'h1f:1'h1];
  assign T15 = T16 == 1'h1;
  assign T16 = queue_io_deq_bits_x[1'h0:1'h0];
  assign T17 = T3 & T18;
  assign T18 = ~ T19;
  assign T19 = T20 ? CreditCon_1_io_almostOut : CreditCon_io_almostOut;
  assign T20 = vcArbiter_io_chosen;
  assign T21 = queue_io_deq_valid | T22;
  assign T22 = 2'h1 <= injQStateMachine_io_currentState;
  assign T23 = T25 | T24;
  assign T24 = 2'h1 <= injQStateMachine_io_currentState;
  assign T25 = CreditCon_io_outCredit & T26;
  assign T26 = T27 == 1'h1;
  assign T27 = queue_io_deq_bits_x[1'h0:1'h0];
  assign T28 = injQStateMachine_io_currentState == 2'h0;
  assign T29 = T31 | T30;
  assign T30 = 2'h1 <= injQStateMachine_io_currentState;
  assign T31 = CreditCon_1_io_outCredit & T32;
  assign T32 = T33 == 1'h1;
  assign T33 = queue_io_deq_bits_x[1'h0:1'h0];
  assign T34 = injQStateMachine_io_currentState == 2'h0;
  assign T35 = T36 & queue_io_deq_valid;
  assign T36 = T37 & T3;
  assign T37 = vcArbiter_io_requests_1_grant & T38;
  assign T38 = injQStateMachine_io_currentState == 2'h2;
  assign T39 = T40 & queue_io_deq_valid;
  assign T40 = T41 & T3;
  assign T41 = vcArbiter_io_requests_0_grant & T42;
  assign T42 = injQStateMachine_io_currentState == 2'h2;
  assign T43 = T0 & queue_io_deq_valid;
  assign io_out_flitValid = T44;
  assign T44 = T45 & queue_io_deq_valid;
  assign T45 = injQStateMachine_io_currentState == 2'h2;
  assign io_out_flit_x = replaceVC_io_newFlit_x;
  assign io_in_credit_grant = creditGen_io_outCredit_grant;
  CreditGen creditGen(
       .io_outCredit_grant( creditGen_io_outCredit_grant ),
       .io_inGrant( T43 )
  );
  CreditCon CreditCon(.clk(clk), .reset(reset),
       .io_inCredit_grant( io_out_credit_0_grant ),
       .io_inConsume( T39 ),
       .io_outCredit( CreditCon_io_outCredit ),
       .io_almostOut( CreditCon_io_almostOut )
  );
  CreditCon CreditCon_1(.clk(clk), .reset(reset),
       .io_inCredit_grant( io_out_credit_1_grant ),
       .io_inConsume( T35 ),
       .io_outCredit( CreditCon_1_io_outCredit ),
       .io_almostOut( CreditCon_1_io_almostOut )
  );
  RRArbiter_0 vcArbiter(.clk(clk), .reset(reset),
       .io_requests_1_releaseLock( T34 ),
       .io_requests_1_grant( vcArbiter_io_requests_1_grant ),
       .io_requests_1_request( T29 ),
       //.io_requests_1_priorityLevel(  )
       .io_requests_0_releaseLock( T28 ),
       .io_requests_0_grant( vcArbiter_io_requests_0_grant ),
       .io_requests_0_request( T23 ),
       //.io_requests_0_priorityLevel(  )
       .io_resource_ready( T21 ),
       .io_resource_valid( vcArbiter_io_resource_valid ),
       .io_chosen( vcArbiter_io_chosen )
  );
  InjectionQStateMgmt injQStateMachine(.clk(clk), .reset(reset),
       .io_inputBufferValid( queue_io_deq_valid ),
       .io_creditsAvailable( T17 ),
       .io_inputIsTail( T8 ),
       .io_vcAllocGranted( vcArbiter_io_resource_valid ),
       .io_currentState( injQStateMachine_io_currentState )
  );
  Queue_0 queue(.clk(clk), .reset(reset),
       //.io_enq_ready(  )
       .io_enq_valid( T5 ),
       .io_enq_bits_x( io_in_flit_x ),
       .io_deq_ready( T0 ),
       .io_deq_valid( queue_io_deq_valid ),
       .io_deq_bits_x( queue_io_deq_bits_x ),
       .io_count( queue_io_count )
  );
  ReplaceVCPort replaceVC(
       .io_oldFlit_x( queue_io_deq_bits_x ),
       .io_newVCPort( vcArbiter_io_chosen ),
       .io_newFlit_x( replaceVC_io_newFlit_x )
  );
endmodule

module Queue_1(input clk, input reset,
    output io_enq_ready,
    input  io_enq_valid,
    input [54:0] io_enq_bits_x,
    input  io_deq_ready,
    output io_deq_valid,
    output[54:0] io_deq_bits_x,
    output[5:0] io_count
);

  wire[5:0] T0;
  wire[4:0] ptr_diff;
  reg [4:0] R1;
  wire[4:0] T16;
  wire[4:0] T2;
  wire[4:0] T3;
  wire do_deq;
  reg [4:0] R4;
  wire[4:0] T17;
  wire[4:0] T5;
  wire[4:0] T6;
  wire do_enq;
  wire T7;
  wire ptr_match;
  reg  maybe_full;
  wire T18;
  wire T8;
  wire T9;
  wire[54:0] T10;
  wire[54:0] T11;
  reg [54:0] ram [31:0];
  wire[54:0] T12;
  wire T13;
  wire empty;
  wire T14;
  wire T15;
  wire full;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    R1 = {1{1'b0}};
    R4 = {1{1'b0}};
    maybe_full = {1{1'b0}};
    for (initvar = 0; initvar < 32; initvar = initvar+1)
      ram[initvar] = {2{1'b0}};
  end
// synthesis translate_on
`endif

  assign io_count = T0;
  assign T0 = {T7, ptr_diff};
  assign ptr_diff = R4 - R1;
  assign T16 = reset ? 5'h0 : T2;
  assign T2 = do_deq ? T3 : R1;
  assign T3 = R1 + 5'h1;
  assign do_deq = io_deq_ready & io_deq_valid;
  assign T17 = reset ? 5'h0 : T5;
  assign T5 = do_enq ? T6 : R4;
  assign T6 = R4 + 5'h1;
  assign do_enq = io_enq_ready & io_enq_valid;
  assign T7 = maybe_full & ptr_match;
  assign ptr_match = R4 == R1;
  assign T18 = reset ? 1'h0 : T8;
  assign T8 = T9 ? do_enq : maybe_full;
  assign T9 = do_enq != do_deq;
  assign io_deq_bits_x = T10;
  assign T10 = T11[6'h36:1'h0];
  assign T11 = ram[R1];
  assign io_deq_valid = T13;
  assign T13 = empty ^ 1'h1;
  assign empty = ptr_match & T14;
  assign T14 = maybe_full ^ 1'h1;
  assign io_enq_ready = T15;
  assign T15 = full ^ 1'h1;
  assign full = ptr_match & maybe_full;

  always @(posedge clk) begin
    if(reset) begin
      R1 <= 5'h0;
    end else if(do_deq) begin
      R1 <= T3;
    end
    if(reset) begin
      R4 <= 5'h0;
    end else if(do_enq) begin
      R4 <= T6;
    end
    if(reset) begin
      maybe_full <= 1'h0;
    end else if(T9) begin
      maybe_full <= do_enq;
    end
    if (do_enq)
      ram[R4] <= io_enq_bits_x;
  end
endmodule

module EjectionChannelQ(input clk, input reset,
    input [54:0] io_in_flit_x,
    input  io_in_flitValid,
    output io_in_credit_1_grant,
    output io_in_credit_0_grant,
    output[54:0] io_out_flit_x,
    output io_out_flitValid,
    input  io_out_credit_grant
);

  wire T0;
  wire T1;
  wire T2;
  wire CreditGen_io_outCredit_grant;
  wire CreditGen_1_io_outCredit_grant;
  wire creditCon_io_outCredit;
  wire queue_io_deq_valid;
  wire[54:0] queue_io_deq_bits_x;


  assign T0 = queue_io_deq_valid & creditCon_io_outCredit;
  assign T1 = creditCon_io_outCredit & queue_io_deq_valid;
  assign T2 = creditCon_io_outCredit & queue_io_deq_valid;
  assign io_out_flitValid = queue_io_deq_valid;
  assign io_out_flit_x = queue_io_deq_bits_x;
  assign io_in_credit_0_grant = CreditGen_io_outCredit_grant;
  assign io_in_credit_1_grant = CreditGen_1_io_outCredit_grant;
  CreditGen CreditGen(
       .io_outCredit_grant( CreditGen_io_outCredit_grant ),
       .io_inGrant( T2 )
  );
  CreditGen CreditGen_1(
       .io_outCredit_grant( CreditGen_1_io_outCredit_grant ),
       .io_inGrant( T1 )
  );
  CreditCon creditCon(.clk(clk), .reset(reset),
       .io_inCredit_grant( io_out_credit_grant ),
       .io_inConsume( T0 ),
       .io_outCredit( creditCon_io_outCredit )
       //.io_almostOut(  )
  );
  Queue_1 queue(.clk(clk), .reset(reset),
       //.io_enq_ready(  )
       .io_enq_valid( io_in_flitValid ),
       .io_enq_bits_x( io_in_flit_x ),
       .io_deq_ready( creditCon_io_outCredit ),
       .io_deq_valid( queue_io_deq_valid ),
       .io_deq_bits_x( queue_io_deq_bits_x )
       //.io_count(  )
  );
endmodule

module FlitToFlit(
    input [54:0] io_packet_x,
    output io_packetReady,
    input  io_packetValid,
    output[54:0] io_flit_x,
    input  io_flitReady,
    output io_flitValid
);



  assign io_flitValid = io_packetValid;
  assign io_flit_x = io_packet_x;
  assign io_packetReady = io_flitReady;
endmodule

module InputPacketInterface(input clk, input reset,
    output io_in_ready,
    input  io_in_valid,
    input [54:0] io_in_bits_x,
    output[54:0] io_out_flit_x,
    output io_out_flitValid,
    input  io_out_credit_grant
);

  wire creditCon_io_outCredit;
  wire packet2Flit_io_packetReady;
  wire[54:0] packet2Flit_io_flit_x;
  wire packet2Flit_io_flitValid;


  assign io_out_flitValid = packet2Flit_io_flitValid;
  assign io_out_flit_x = packet2Flit_io_flit_x;
  assign io_in_ready = packet2Flit_io_packetReady;
  CreditCon creditCon(.clk(clk), .reset(reset),
       .io_inCredit_grant( io_out_credit_grant ),
       .io_inConsume( packet2Flit_io_flitValid ),
       .io_outCredit( creditCon_io_outCredit )
       //.io_almostOut(  )
  );
  FlitToFlit packet2Flit(
       .io_packet_x( io_in_bits_x ),
       .io_packetReady( packet2Flit_io_packetReady ),
       .io_packetValid( io_in_valid ),
       .io_flit_x( packet2Flit_io_flit_x ),
       .io_flitReady( creditCon_io_outCredit ),
       .io_flitValid( packet2Flit_io_flitValid )
  );
endmodule

module My_Mesh(input clk, input reset,
    input [54:0] io_ports_2_in_packet_x,
    output io_ports_2_in_packetReady,
    input  io_ports_2_in_packetValid,
    output[54:0] io_ports_2_out_flit_x,
    output io_ports_2_out_flitValid,
    input  io_ports_2_out_credit_grant,
    input [54:0] io_ports_1_in_packet_x,
    output io_ports_1_in_packetReady,
    input  io_ports_1_in_packetValid,
    output[54:0] io_ports_1_out_flit_x,
    output io_ports_1_out_flitValid,
    input  io_ports_1_out_credit_grant,
    input [54:0] io_ports_0_in_packet_x,
    output io_ports_0_in_packetReady,
    input  io_ports_0_in_packetValid,
    output[54:0] io_ports_0_out_flit_x,
    output io_ports_0_out_flitValid,
    input  io_ports_0_out_credit_grant,
    input  io_bypass_2,
    input  io_bypass_1,
    input  io_bypass_0,
    output[15:0] io_cyclesRouterBusy_2,
    output[15:0] io_cyclesRouterBusy_1,
    output[15:0] io_cyclesRouterBusy_0,
    output[15:0] io_cyclesChannelBusy_14,
    output[15:0] io_cyclesChannelBusy_13,
    output[15:0] io_cyclesChannelBusy_12,
    output[15:0] io_cyclesChannelBusy_11,
    output[15:0] io_cyclesChannelBusy_10,
    output[15:0] io_cyclesChannelBusy_9,
    output[15:0] io_cyclesChannelBusy_8,
    output[15:0] io_cyclesChannelBusy_7,
    output[15:0] io_cyclesChannelBusy_6,
    output[15:0] io_cyclesChannelBusy_5,
    output[15:0] io_cyclesChannelBusy_4,
    output[15:0] io_cyclesChannelBusy_3,
    output[15:0] io_cyclesChannelBusy_2,
    output[15:0] io_cyclesChannelBusy_1,
    output[15:0] io_cyclesChannelBusy_0
);

  wire EjectionChannelQ_io_in_credit_1_grant;
  wire EjectionChannelQ_io_in_credit_0_grant;
  wire[54:0] EjectionChannelQ_io_out_flit_x;
  wire EjectionChannelQ_io_out_flitValid;
  wire InputPacketInterface_io_in_ready;
  wire[54:0] InputPacketInterface_io_out_flit_x;
  wire InputPacketInterface_io_out_flitValid;
  wire EjectionChannelQ_1_io_in_credit_1_grant;
  wire EjectionChannelQ_1_io_in_credit_0_grant;
  wire[54:0] EjectionChannelQ_1_io_out_flit_x;
  wire EjectionChannelQ_1_io_out_flitValid;
  wire InputPacketInterface_1_io_in_ready;
  wire[54:0] InputPacketInterface_1_io_out_flit_x;
  wire InputPacketInterface_1_io_out_flitValid;
  wire EjectionChannelQ_2_io_in_credit_1_grant;
  wire EjectionChannelQ_2_io_in_credit_0_grant;
  wire[54:0] EjectionChannelQ_2_io_out_flit_x;
  wire EjectionChannelQ_2_io_out_flitValid;
  wire InputPacketInterface_2_io_in_ready;
  wire[54:0] InputPacketInterface_2_io_out_flit_x;
  wire InputPacketInterface_2_io_out_flitValid;
  wire InjectionChannelQ_io_in_credit_grant;
  wire[54:0] InjectionChannelQ_io_out_flit_x;
  wire InjectionChannelQ_io_out_flitValid;
  wire InjectionChannelQ_1_io_in_credit_grant;
  wire[54:0] InjectionChannelQ_1_io_out_flit_x;
  wire InjectionChannelQ_1_io_out_flitValid;
  wire InjectionChannelQ_2_io_in_credit_grant;
  wire[54:0] InjectionChannelQ_2_io_out_flit_x;
  wire InjectionChannelQ_2_io_out_flitValid;
  wire VCCMesh_io_inChannels_2_credit_1_grant;
  wire VCCMesh_io_inChannels_2_credit_0_grant;
  wire VCCMesh_io_inChannels_1_credit_1_grant;
  wire VCCMesh_io_inChannels_1_credit_0_grant;
  wire VCCMesh_io_inChannels_0_credit_1_grant;
  wire VCCMesh_io_inChannels_0_credit_0_grant;
  wire[54:0] VCCMesh_io_outChannels_2_flit_x;
  wire VCCMesh_io_outChannels_2_flitValid;
  wire[54:0] VCCMesh_io_outChannels_1_flit_x;
  wire VCCMesh_io_outChannels_1_flitValid;
  wire[54:0] VCCMesh_io_outChannels_0_flit_x;
  wire VCCMesh_io_outChannels_0_flitValid;
  wire[15:0] VCCMesh_io_cyclesRouterBusy_2;
  wire[15:0] VCCMesh_io_cyclesRouterBusy_1;
  wire[15:0] VCCMesh_io_cyclesRouterBusy_0;
  wire[15:0] VCCMesh_io_cyclesChannelBusy_14;
  wire[15:0] VCCMesh_io_cyclesChannelBusy_13;
  wire[15:0] VCCMesh_io_cyclesChannelBusy_12;
  wire[15:0] VCCMesh_io_cyclesChannelBusy_11;
  wire[15:0] VCCMesh_io_cyclesChannelBusy_10;
  wire[15:0] VCCMesh_io_cyclesChannelBusy_9;
  wire[15:0] VCCMesh_io_cyclesChannelBusy_8;
  wire[15:0] VCCMesh_io_cyclesChannelBusy_7;
  wire[15:0] VCCMesh_io_cyclesChannelBusy_6;
  wire[15:0] VCCMesh_io_cyclesChannelBusy_5;
  wire[15:0] VCCMesh_io_cyclesChannelBusy_4;
  wire[15:0] VCCMesh_io_cyclesChannelBusy_3;
  wire[15:0] VCCMesh_io_cyclesChannelBusy_2;
  wire[15:0] VCCMesh_io_cyclesChannelBusy_1;
  wire[15:0] VCCMesh_io_cyclesChannelBusy_0;


  assign io_cyclesChannelBusy_0 = VCCMesh_io_cyclesChannelBusy_0;
  assign io_cyclesChannelBusy_1 = VCCMesh_io_cyclesChannelBusy_1;
  assign io_cyclesChannelBusy_2 = VCCMesh_io_cyclesChannelBusy_2;
  assign io_cyclesChannelBusy_3 = VCCMesh_io_cyclesChannelBusy_3;
  assign io_cyclesChannelBusy_4 = VCCMesh_io_cyclesChannelBusy_4;
  assign io_cyclesChannelBusy_5 = VCCMesh_io_cyclesChannelBusy_5;
  assign io_cyclesChannelBusy_6 = VCCMesh_io_cyclesChannelBusy_6;
  assign io_cyclesChannelBusy_7 = VCCMesh_io_cyclesChannelBusy_7;
  assign io_cyclesChannelBusy_8 = VCCMesh_io_cyclesChannelBusy_8;
  assign io_cyclesChannelBusy_9 = VCCMesh_io_cyclesChannelBusy_9;
  assign io_cyclesChannelBusy_10 = VCCMesh_io_cyclesChannelBusy_10;
  assign io_cyclesChannelBusy_11 = VCCMesh_io_cyclesChannelBusy_11;
  assign io_cyclesChannelBusy_12 = VCCMesh_io_cyclesChannelBusy_12;
  assign io_cyclesChannelBusy_13 = VCCMesh_io_cyclesChannelBusy_13;
  assign io_cyclesChannelBusy_14 = VCCMesh_io_cyclesChannelBusy_14;
  assign io_cyclesRouterBusy_0 = VCCMesh_io_cyclesRouterBusy_0;
  assign io_cyclesRouterBusy_1 = VCCMesh_io_cyclesRouterBusy_1;
  assign io_cyclesRouterBusy_2 = VCCMesh_io_cyclesRouterBusy_2;
  assign io_ports_0_out_flitValid = EjectionChannelQ_io_out_flitValid;
  assign io_ports_0_out_flit_x = EjectionChannelQ_io_out_flit_x;
  assign io_ports_0_in_packetReady = InputPacketInterface_io_in_ready;
  assign io_ports_1_out_flitValid = EjectionChannelQ_1_io_out_flitValid;
  assign io_ports_1_out_flit_x = EjectionChannelQ_1_io_out_flit_x;
  assign io_ports_1_in_packetReady = InputPacketInterface_1_io_in_ready;
  assign io_ports_2_out_flitValid = EjectionChannelQ_2_io_out_flitValid;
  assign io_ports_2_out_flit_x = EjectionChannelQ_2_io_out_flit_x;
  assign io_ports_2_in_packetReady = InputPacketInterface_2_io_in_ready;
  VCCMesh VCCMesh(.clk(clk), .reset(reset),
       .io_inChannels_2_flit_x( InjectionChannelQ_2_io_out_flit_x ),
       .io_inChannels_2_flitValid( InjectionChannelQ_2_io_out_flitValid ),
       .io_inChannels_2_credit_1_grant( VCCMesh_io_inChannels_2_credit_1_grant ),
       .io_inChannels_2_credit_0_grant( VCCMesh_io_inChannels_2_credit_0_grant ),
       .io_inChannels_1_flit_x( InjectionChannelQ_1_io_out_flit_x ),
       .io_inChannels_1_flitValid( InjectionChannelQ_1_io_out_flitValid ),
       .io_inChannels_1_credit_1_grant( VCCMesh_io_inChannels_1_credit_1_grant ),
       .io_inChannels_1_credit_0_grant( VCCMesh_io_inChannels_1_credit_0_grant ),
       .io_inChannels_0_flit_x( InjectionChannelQ_io_out_flit_x ),
       .io_inChannels_0_flitValid( InjectionChannelQ_io_out_flitValid ),
       .io_inChannels_0_credit_1_grant( VCCMesh_io_inChannels_0_credit_1_grant ),
       .io_inChannels_0_credit_0_grant( VCCMesh_io_inChannels_0_credit_0_grant ),
       .io_outChannels_2_flit_x( VCCMesh_io_outChannels_2_flit_x ),
       .io_outChannels_2_flitValid( VCCMesh_io_outChannels_2_flitValid ),
       .io_outChannels_2_credit_1_grant( EjectionChannelQ_2_io_in_credit_1_grant ),
       .io_outChannels_2_credit_0_grant( EjectionChannelQ_2_io_in_credit_0_grant ),
       .io_outChannels_1_flit_x( VCCMesh_io_outChannels_1_flit_x ),
       .io_outChannels_1_flitValid( VCCMesh_io_outChannels_1_flitValid ),
       .io_outChannels_1_credit_1_grant( EjectionChannelQ_1_io_in_credit_1_grant ),
       .io_outChannels_1_credit_0_grant( EjectionChannelQ_1_io_in_credit_0_grant ),
       .io_outChannels_0_flit_x( VCCMesh_io_outChannels_0_flit_x ),
       .io_outChannels_0_flitValid( VCCMesh_io_outChannels_0_flitValid ),
       .io_outChannels_0_credit_1_grant( EjectionChannelQ_io_in_credit_1_grant ),
       .io_outChannels_0_credit_0_grant( EjectionChannelQ_io_in_credit_0_grant ),
       //.io_cyclesRouterBusy_127(  )
       //.io_cyclesRouterBusy_126(  )
       //.io_cyclesRouterBusy_125(  )
       //.io_cyclesRouterBusy_124(  )
       //.io_cyclesRouterBusy_123(  )
       //.io_cyclesRouterBusy_122(  )
       //.io_cyclesRouterBusy_121(  )
       //.io_cyclesRouterBusy_120(  )
       //.io_cyclesRouterBusy_119(  )
       //.io_cyclesRouterBusy_118(  )
       //.io_cyclesRouterBusy_117(  )
       //.io_cyclesRouterBusy_116(  )
       //.io_cyclesRouterBusy_115(  )
       //.io_cyclesRouterBusy_114(  )
       //.io_cyclesRouterBusy_113(  )
       //.io_cyclesRouterBusy_112(  )
       //.io_cyclesRouterBusy_111(  )
       //.io_cyclesRouterBusy_110(  )
       //.io_cyclesRouterBusy_109(  )
       //.io_cyclesRouterBusy_108(  )
       //.io_cyclesRouterBusy_107(  )
       //.io_cyclesRouterBusy_106(  )
       //.io_cyclesRouterBusy_105(  )
       //.io_cyclesRouterBusy_104(  )
       //.io_cyclesRouterBusy_103(  )
       //.io_cyclesRouterBusy_102(  )
       //.io_cyclesRouterBusy_101(  )
       //.io_cyclesRouterBusy_100(  )
       //.io_cyclesRouterBusy_99(  )
       //.io_cyclesRouterBusy_98(  )
       //.io_cyclesRouterBusy_97(  )
       //.io_cyclesRouterBusy_96(  )
       //.io_cyclesRouterBusy_95(  )
       //.io_cyclesRouterBusy_94(  )
       //.io_cyclesRouterBusy_93(  )
       //.io_cyclesRouterBusy_92(  )
       //.io_cyclesRouterBusy_91(  )
       //.io_cyclesRouterBusy_90(  )
       //.io_cyclesRouterBusy_89(  )
       //.io_cyclesRouterBusy_88(  )
       //.io_cyclesRouterBusy_87(  )
       //.io_cyclesRouterBusy_86(  )
       //.io_cyclesRouterBusy_85(  )
       //.io_cyclesRouterBusy_84(  )
       //.io_cyclesRouterBusy_83(  )
       //.io_cyclesRouterBusy_82(  )
       //.io_cyclesRouterBusy_81(  )
       //.io_cyclesRouterBusy_80(  )
       //.io_cyclesRouterBusy_79(  )
       //.io_cyclesRouterBusy_78(  )
       //.io_cyclesRouterBusy_77(  )
       //.io_cyclesRouterBusy_76(  )
       //.io_cyclesRouterBusy_75(  )
       //.io_cyclesRouterBusy_74(  )
       //.io_cyclesRouterBusy_73(  )
       //.io_cyclesRouterBusy_72(  )
       //.io_cyclesRouterBusy_71(  )
       //.io_cyclesRouterBusy_70(  )
       //.io_cyclesRouterBusy_69(  )
       //.io_cyclesRouterBusy_68(  )
       //.io_cyclesRouterBusy_67(  )
       //.io_cyclesRouterBusy_66(  )
       //.io_cyclesRouterBusy_65(  )
       //.io_cyclesRouterBusy_64(  )
       //.io_cyclesRouterBusy_63(  )
       //.io_cyclesRouterBusy_62(  )
       //.io_cyclesRouterBusy_61(  )
       //.io_cyclesRouterBusy_60(  )
       //.io_cyclesRouterBusy_59(  )
       //.io_cyclesRouterBusy_58(  )
       //.io_cyclesRouterBusy_57(  )
       //.io_cyclesRouterBusy_56(  )
       //.io_cyclesRouterBusy_55(  )
       //.io_cyclesRouterBusy_54(  )
       //.io_cyclesRouterBusy_53(  )
       //.io_cyclesRouterBusy_52(  )
       //.io_cyclesRouterBusy_51(  )
       //.io_cyclesRouterBusy_50(  )
       //.io_cyclesRouterBusy_49(  )
       //.io_cyclesRouterBusy_48(  )
       //.io_cyclesRouterBusy_47(  )
       //.io_cyclesRouterBusy_46(  )
       //.io_cyclesRouterBusy_45(  )
       //.io_cyclesRouterBusy_44(  )
       //.io_cyclesRouterBusy_43(  )
       //.io_cyclesRouterBusy_42(  )
       //.io_cyclesRouterBusy_41(  )
       //.io_cyclesRouterBusy_40(  )
       //.io_cyclesRouterBusy_39(  )
       //.io_cyclesRouterBusy_38(  )
       //.io_cyclesRouterBusy_37(  )
       //.io_cyclesRouterBusy_36(  )
       //.io_cyclesRouterBusy_35(  )
       //.io_cyclesRouterBusy_34(  )
       //.io_cyclesRouterBusy_33(  )
       //.io_cyclesRouterBusy_32(  )
       //.io_cyclesRouterBusy_31(  )
       //.io_cyclesRouterBusy_30(  )
       //.io_cyclesRouterBusy_29(  )
       //.io_cyclesRouterBusy_28(  )
       //.io_cyclesRouterBusy_27(  )
       //.io_cyclesRouterBusy_26(  )
       //.io_cyclesRouterBusy_25(  )
       //.io_cyclesRouterBusy_24(  )
       //.io_cyclesRouterBusy_23(  )
       //.io_cyclesRouterBusy_22(  )
       //.io_cyclesRouterBusy_21(  )
       //.io_cyclesRouterBusy_20(  )
       //.io_cyclesRouterBusy_19(  )
       //.io_cyclesRouterBusy_18(  )
       //.io_cyclesRouterBusy_17(  )
       //.io_cyclesRouterBusy_16(  )
       //.io_cyclesRouterBusy_15(  )
       //.io_cyclesRouterBusy_14(  )
       //.io_cyclesRouterBusy_13(  )
       //.io_cyclesRouterBusy_12(  )
       //.io_cyclesRouterBusy_11(  )
       //.io_cyclesRouterBusy_10(  )
       //.io_cyclesRouterBusy_9(  )
       //.io_cyclesRouterBusy_8(  )
       //.io_cyclesRouterBusy_7(  )
       //.io_cyclesRouterBusy_6(  )
       //.io_cyclesRouterBusy_5(  )
       //.io_cyclesRouterBusy_4(  )
       //.io_cyclesRouterBusy_3(  )
       .io_cyclesRouterBusy_2( VCCMesh_io_cyclesRouterBusy_2 ),
       .io_cyclesRouterBusy_1( VCCMesh_io_cyclesRouterBusy_1 ),
       .io_cyclesRouterBusy_0( VCCMesh_io_cyclesRouterBusy_0 ),
       //.io_cyclesChannelBusy_639(  )
       //.io_cyclesChannelBusy_638(  )
       //.io_cyclesChannelBusy_637(  )
       //.io_cyclesChannelBusy_636(  )
       //.io_cyclesChannelBusy_635(  )
       //.io_cyclesChannelBusy_634(  )
       //.io_cyclesChannelBusy_633(  )
       //.io_cyclesChannelBusy_632(  )
       //.io_cyclesChannelBusy_631(  )
       //.io_cyclesChannelBusy_630(  )
       //.io_cyclesChannelBusy_629(  )
       //.io_cyclesChannelBusy_628(  )
       //.io_cyclesChannelBusy_627(  )
       //.io_cyclesChannelBusy_626(  )
       //.io_cyclesChannelBusy_625(  )
       //.io_cyclesChannelBusy_624(  )
       //.io_cyclesChannelBusy_623(  )
       //.io_cyclesChannelBusy_622(  )
       //.io_cyclesChannelBusy_621(  )
       //.io_cyclesChannelBusy_620(  )
       //.io_cyclesChannelBusy_619(  )
       //.io_cyclesChannelBusy_618(  )
       //.io_cyclesChannelBusy_617(  )
       //.io_cyclesChannelBusy_616(  )
       //.io_cyclesChannelBusy_615(  )
       //.io_cyclesChannelBusy_614(  )
       //.io_cyclesChannelBusy_613(  )
       //.io_cyclesChannelBusy_612(  )
       //.io_cyclesChannelBusy_611(  )
       //.io_cyclesChannelBusy_610(  )
       //.io_cyclesChannelBusy_609(  )
       //.io_cyclesChannelBusy_608(  )
       //.io_cyclesChannelBusy_607(  )
       //.io_cyclesChannelBusy_606(  )
       //.io_cyclesChannelBusy_605(  )
       //.io_cyclesChannelBusy_604(  )
       //.io_cyclesChannelBusy_603(  )
       //.io_cyclesChannelBusy_602(  )
       //.io_cyclesChannelBusy_601(  )
       //.io_cyclesChannelBusy_600(  )
       //.io_cyclesChannelBusy_599(  )
       //.io_cyclesChannelBusy_598(  )
       //.io_cyclesChannelBusy_597(  )
       //.io_cyclesChannelBusy_596(  )
       //.io_cyclesChannelBusy_595(  )
       //.io_cyclesChannelBusy_594(  )
       //.io_cyclesChannelBusy_593(  )
       //.io_cyclesChannelBusy_592(  )
       //.io_cyclesChannelBusy_591(  )
       //.io_cyclesChannelBusy_590(  )
       //.io_cyclesChannelBusy_589(  )
       //.io_cyclesChannelBusy_588(  )
       //.io_cyclesChannelBusy_587(  )
       //.io_cyclesChannelBusy_586(  )
       //.io_cyclesChannelBusy_585(  )
       //.io_cyclesChannelBusy_584(  )
       //.io_cyclesChannelBusy_583(  )
       //.io_cyclesChannelBusy_582(  )
       //.io_cyclesChannelBusy_581(  )
       //.io_cyclesChannelBusy_580(  )
       //.io_cyclesChannelBusy_579(  )
       //.io_cyclesChannelBusy_578(  )
       //.io_cyclesChannelBusy_577(  )
       //.io_cyclesChannelBusy_576(  )
       //.io_cyclesChannelBusy_575(  )
       //.io_cyclesChannelBusy_574(  )
       //.io_cyclesChannelBusy_573(  )
       //.io_cyclesChannelBusy_572(  )
       //.io_cyclesChannelBusy_571(  )
       //.io_cyclesChannelBusy_570(  )
       //.io_cyclesChannelBusy_569(  )
       //.io_cyclesChannelBusy_568(  )
       //.io_cyclesChannelBusy_567(  )
       //.io_cyclesChannelBusy_566(  )
       //.io_cyclesChannelBusy_565(  )
       //.io_cyclesChannelBusy_564(  )
       //.io_cyclesChannelBusy_563(  )
       //.io_cyclesChannelBusy_562(  )
       //.io_cyclesChannelBusy_561(  )
       //.io_cyclesChannelBusy_560(  )
       //.io_cyclesChannelBusy_559(  )
       //.io_cyclesChannelBusy_558(  )
       //.io_cyclesChannelBusy_557(  )
       //.io_cyclesChannelBusy_556(  )
       //.io_cyclesChannelBusy_555(  )
       //.io_cyclesChannelBusy_554(  )
       //.io_cyclesChannelBusy_553(  )
       //.io_cyclesChannelBusy_552(  )
       //.io_cyclesChannelBusy_551(  )
       //.io_cyclesChannelBusy_550(  )
       //.io_cyclesChannelBusy_549(  )
       //.io_cyclesChannelBusy_548(  )
       //.io_cyclesChannelBusy_547(  )
       //.io_cyclesChannelBusy_546(  )
       //.io_cyclesChannelBusy_545(  )
       //.io_cyclesChannelBusy_544(  )
       //.io_cyclesChannelBusy_543(  )
       //.io_cyclesChannelBusy_542(  )
       //.io_cyclesChannelBusy_541(  )
       //.io_cyclesChannelBusy_540(  )
       //.io_cyclesChannelBusy_539(  )
       //.io_cyclesChannelBusy_538(  )
       //.io_cyclesChannelBusy_537(  )
       //.io_cyclesChannelBusy_536(  )
       //.io_cyclesChannelBusy_535(  )
       //.io_cyclesChannelBusy_534(  )
       //.io_cyclesChannelBusy_533(  )
       //.io_cyclesChannelBusy_532(  )
       //.io_cyclesChannelBusy_531(  )
       //.io_cyclesChannelBusy_530(  )
       //.io_cyclesChannelBusy_529(  )
       //.io_cyclesChannelBusy_528(  )
       //.io_cyclesChannelBusy_527(  )
       //.io_cyclesChannelBusy_526(  )
       //.io_cyclesChannelBusy_525(  )
       //.io_cyclesChannelBusy_524(  )
       //.io_cyclesChannelBusy_523(  )
       //.io_cyclesChannelBusy_522(  )
       //.io_cyclesChannelBusy_521(  )
       //.io_cyclesChannelBusy_520(  )
       //.io_cyclesChannelBusy_519(  )
       //.io_cyclesChannelBusy_518(  )
       //.io_cyclesChannelBusy_517(  )
       //.io_cyclesChannelBusy_516(  )
       //.io_cyclesChannelBusy_515(  )
       //.io_cyclesChannelBusy_514(  )
       //.io_cyclesChannelBusy_513(  )
       //.io_cyclesChannelBusy_512(  )
       //.io_cyclesChannelBusy_511(  )
       //.io_cyclesChannelBusy_510(  )
       //.io_cyclesChannelBusy_509(  )
       //.io_cyclesChannelBusy_508(  )
       //.io_cyclesChannelBusy_507(  )
       //.io_cyclesChannelBusy_506(  )
       //.io_cyclesChannelBusy_505(  )
       //.io_cyclesChannelBusy_504(  )
       //.io_cyclesChannelBusy_503(  )
       //.io_cyclesChannelBusy_502(  )
       //.io_cyclesChannelBusy_501(  )
       //.io_cyclesChannelBusy_500(  )
       //.io_cyclesChannelBusy_499(  )
       //.io_cyclesChannelBusy_498(  )
       //.io_cyclesChannelBusy_497(  )
       //.io_cyclesChannelBusy_496(  )
       //.io_cyclesChannelBusy_495(  )
       //.io_cyclesChannelBusy_494(  )
       //.io_cyclesChannelBusy_493(  )
       //.io_cyclesChannelBusy_492(  )
       //.io_cyclesChannelBusy_491(  )
       //.io_cyclesChannelBusy_490(  )
       //.io_cyclesChannelBusy_489(  )
       //.io_cyclesChannelBusy_488(  )
       //.io_cyclesChannelBusy_487(  )
       //.io_cyclesChannelBusy_486(  )
       //.io_cyclesChannelBusy_485(  )
       //.io_cyclesChannelBusy_484(  )
       //.io_cyclesChannelBusy_483(  )
       //.io_cyclesChannelBusy_482(  )
       //.io_cyclesChannelBusy_481(  )
       //.io_cyclesChannelBusy_480(  )
       //.io_cyclesChannelBusy_479(  )
       //.io_cyclesChannelBusy_478(  )
       //.io_cyclesChannelBusy_477(  )
       //.io_cyclesChannelBusy_476(  )
       //.io_cyclesChannelBusy_475(  )
       //.io_cyclesChannelBusy_474(  )
       //.io_cyclesChannelBusy_473(  )
       //.io_cyclesChannelBusy_472(  )
       //.io_cyclesChannelBusy_471(  )
       //.io_cyclesChannelBusy_470(  )
       //.io_cyclesChannelBusy_469(  )
       //.io_cyclesChannelBusy_468(  )
       //.io_cyclesChannelBusy_467(  )
       //.io_cyclesChannelBusy_466(  )
       //.io_cyclesChannelBusy_465(  )
       //.io_cyclesChannelBusy_464(  )
       //.io_cyclesChannelBusy_463(  )
       //.io_cyclesChannelBusy_462(  )
       //.io_cyclesChannelBusy_461(  )
       //.io_cyclesChannelBusy_460(  )
       //.io_cyclesChannelBusy_459(  )
       //.io_cyclesChannelBusy_458(  )
       //.io_cyclesChannelBusy_457(  )
       //.io_cyclesChannelBusy_456(  )
       //.io_cyclesChannelBusy_455(  )
       //.io_cyclesChannelBusy_454(  )
       //.io_cyclesChannelBusy_453(  )
       //.io_cyclesChannelBusy_452(  )
       //.io_cyclesChannelBusy_451(  )
       //.io_cyclesChannelBusy_450(  )
       //.io_cyclesChannelBusy_449(  )
       //.io_cyclesChannelBusy_448(  )
       //.io_cyclesChannelBusy_447(  )
       //.io_cyclesChannelBusy_446(  )
       //.io_cyclesChannelBusy_445(  )
       //.io_cyclesChannelBusy_444(  )
       //.io_cyclesChannelBusy_443(  )
       //.io_cyclesChannelBusy_442(  )
       //.io_cyclesChannelBusy_441(  )
       //.io_cyclesChannelBusy_440(  )
       //.io_cyclesChannelBusy_439(  )
       //.io_cyclesChannelBusy_438(  )
       //.io_cyclesChannelBusy_437(  )
       //.io_cyclesChannelBusy_436(  )
       //.io_cyclesChannelBusy_435(  )
       //.io_cyclesChannelBusy_434(  )
       //.io_cyclesChannelBusy_433(  )
       //.io_cyclesChannelBusy_432(  )
       //.io_cyclesChannelBusy_431(  )
       //.io_cyclesChannelBusy_430(  )
       //.io_cyclesChannelBusy_429(  )
       //.io_cyclesChannelBusy_428(  )
       //.io_cyclesChannelBusy_427(  )
       //.io_cyclesChannelBusy_426(  )
       //.io_cyclesChannelBusy_425(  )
       //.io_cyclesChannelBusy_424(  )
       //.io_cyclesChannelBusy_423(  )
       //.io_cyclesChannelBusy_422(  )
       //.io_cyclesChannelBusy_421(  )
       //.io_cyclesChannelBusy_420(  )
       //.io_cyclesChannelBusy_419(  )
       //.io_cyclesChannelBusy_418(  )
       //.io_cyclesChannelBusy_417(  )
       //.io_cyclesChannelBusy_416(  )
       //.io_cyclesChannelBusy_415(  )
       //.io_cyclesChannelBusy_414(  )
       //.io_cyclesChannelBusy_413(  )
       //.io_cyclesChannelBusy_412(  )
       //.io_cyclesChannelBusy_411(  )
       //.io_cyclesChannelBusy_410(  )
       //.io_cyclesChannelBusy_409(  )
       //.io_cyclesChannelBusy_408(  )
       //.io_cyclesChannelBusy_407(  )
       //.io_cyclesChannelBusy_406(  )
       //.io_cyclesChannelBusy_405(  )
       //.io_cyclesChannelBusy_404(  )
       //.io_cyclesChannelBusy_403(  )
       //.io_cyclesChannelBusy_402(  )
       //.io_cyclesChannelBusy_401(  )
       //.io_cyclesChannelBusy_400(  )
       //.io_cyclesChannelBusy_399(  )
       //.io_cyclesChannelBusy_398(  )
       //.io_cyclesChannelBusy_397(  )
       //.io_cyclesChannelBusy_396(  )
       //.io_cyclesChannelBusy_395(  )
       //.io_cyclesChannelBusy_394(  )
       //.io_cyclesChannelBusy_393(  )
       //.io_cyclesChannelBusy_392(  )
       //.io_cyclesChannelBusy_391(  )
       //.io_cyclesChannelBusy_390(  )
       //.io_cyclesChannelBusy_389(  )
       //.io_cyclesChannelBusy_388(  )
       //.io_cyclesChannelBusy_387(  )
       //.io_cyclesChannelBusy_386(  )
       //.io_cyclesChannelBusy_385(  )
       //.io_cyclesChannelBusy_384(  )
       //.io_cyclesChannelBusy_383(  )
       //.io_cyclesChannelBusy_382(  )
       //.io_cyclesChannelBusy_381(  )
       //.io_cyclesChannelBusy_380(  )
       //.io_cyclesChannelBusy_379(  )
       //.io_cyclesChannelBusy_378(  )
       //.io_cyclesChannelBusy_377(  )
       //.io_cyclesChannelBusy_376(  )
       //.io_cyclesChannelBusy_375(  )
       //.io_cyclesChannelBusy_374(  )
       //.io_cyclesChannelBusy_373(  )
       //.io_cyclesChannelBusy_372(  )
       //.io_cyclesChannelBusy_371(  )
       //.io_cyclesChannelBusy_370(  )
       //.io_cyclesChannelBusy_369(  )
       //.io_cyclesChannelBusy_368(  )
       //.io_cyclesChannelBusy_367(  )
       //.io_cyclesChannelBusy_366(  )
       //.io_cyclesChannelBusy_365(  )
       //.io_cyclesChannelBusy_364(  )
       //.io_cyclesChannelBusy_363(  )
       //.io_cyclesChannelBusy_362(  )
       //.io_cyclesChannelBusy_361(  )
       //.io_cyclesChannelBusy_360(  )
       //.io_cyclesChannelBusy_359(  )
       //.io_cyclesChannelBusy_358(  )
       //.io_cyclesChannelBusy_357(  )
       //.io_cyclesChannelBusy_356(  )
       //.io_cyclesChannelBusy_355(  )
       //.io_cyclesChannelBusy_354(  )
       //.io_cyclesChannelBusy_353(  )
       //.io_cyclesChannelBusy_352(  )
       //.io_cyclesChannelBusy_351(  )
       //.io_cyclesChannelBusy_350(  )
       //.io_cyclesChannelBusy_349(  )
       //.io_cyclesChannelBusy_348(  )
       //.io_cyclesChannelBusy_347(  )
       //.io_cyclesChannelBusy_346(  )
       //.io_cyclesChannelBusy_345(  )
       //.io_cyclesChannelBusy_344(  )
       //.io_cyclesChannelBusy_343(  )
       //.io_cyclesChannelBusy_342(  )
       //.io_cyclesChannelBusy_341(  )
       //.io_cyclesChannelBusy_340(  )
       //.io_cyclesChannelBusy_339(  )
       //.io_cyclesChannelBusy_338(  )
       //.io_cyclesChannelBusy_337(  )
       //.io_cyclesChannelBusy_336(  )
       //.io_cyclesChannelBusy_335(  )
       //.io_cyclesChannelBusy_334(  )
       //.io_cyclesChannelBusy_333(  )
       //.io_cyclesChannelBusy_332(  )
       //.io_cyclesChannelBusy_331(  )
       //.io_cyclesChannelBusy_330(  )
       //.io_cyclesChannelBusy_329(  )
       //.io_cyclesChannelBusy_328(  )
       //.io_cyclesChannelBusy_327(  )
       //.io_cyclesChannelBusy_326(  )
       //.io_cyclesChannelBusy_325(  )
       //.io_cyclesChannelBusy_324(  )
       //.io_cyclesChannelBusy_323(  )
       //.io_cyclesChannelBusy_322(  )
       //.io_cyclesChannelBusy_321(  )
       //.io_cyclesChannelBusy_320(  )
       //.io_cyclesChannelBusy_319(  )
       //.io_cyclesChannelBusy_318(  )
       //.io_cyclesChannelBusy_317(  )
       //.io_cyclesChannelBusy_316(  )
       //.io_cyclesChannelBusy_315(  )
       //.io_cyclesChannelBusy_314(  )
       //.io_cyclesChannelBusy_313(  )
       //.io_cyclesChannelBusy_312(  )
       //.io_cyclesChannelBusy_311(  )
       //.io_cyclesChannelBusy_310(  )
       //.io_cyclesChannelBusy_309(  )
       //.io_cyclesChannelBusy_308(  )
       //.io_cyclesChannelBusy_307(  )
       //.io_cyclesChannelBusy_306(  )
       //.io_cyclesChannelBusy_305(  )
       //.io_cyclesChannelBusy_304(  )
       //.io_cyclesChannelBusy_303(  )
       //.io_cyclesChannelBusy_302(  )
       //.io_cyclesChannelBusy_301(  )
       //.io_cyclesChannelBusy_300(  )
       //.io_cyclesChannelBusy_299(  )
       //.io_cyclesChannelBusy_298(  )
       //.io_cyclesChannelBusy_297(  )
       //.io_cyclesChannelBusy_296(  )
       //.io_cyclesChannelBusy_295(  )
       //.io_cyclesChannelBusy_294(  )
       //.io_cyclesChannelBusy_293(  )
       //.io_cyclesChannelBusy_292(  )
       //.io_cyclesChannelBusy_291(  )
       //.io_cyclesChannelBusy_290(  )
       //.io_cyclesChannelBusy_289(  )
       //.io_cyclesChannelBusy_288(  )
       //.io_cyclesChannelBusy_287(  )
       //.io_cyclesChannelBusy_286(  )
       //.io_cyclesChannelBusy_285(  )
       //.io_cyclesChannelBusy_284(  )
       //.io_cyclesChannelBusy_283(  )
       //.io_cyclesChannelBusy_282(  )
       //.io_cyclesChannelBusy_281(  )
       //.io_cyclesChannelBusy_280(  )
       //.io_cyclesChannelBusy_279(  )
       //.io_cyclesChannelBusy_278(  )
       //.io_cyclesChannelBusy_277(  )
       //.io_cyclesChannelBusy_276(  )
       //.io_cyclesChannelBusy_275(  )
       //.io_cyclesChannelBusy_274(  )
       //.io_cyclesChannelBusy_273(  )
       //.io_cyclesChannelBusy_272(  )
       //.io_cyclesChannelBusy_271(  )
       //.io_cyclesChannelBusy_270(  )
       //.io_cyclesChannelBusy_269(  )
       //.io_cyclesChannelBusy_268(  )
       //.io_cyclesChannelBusy_267(  )
       //.io_cyclesChannelBusy_266(  )
       //.io_cyclesChannelBusy_265(  )
       //.io_cyclesChannelBusy_264(  )
       //.io_cyclesChannelBusy_263(  )
       //.io_cyclesChannelBusy_262(  )
       //.io_cyclesChannelBusy_261(  )
       //.io_cyclesChannelBusy_260(  )
       //.io_cyclesChannelBusy_259(  )
       //.io_cyclesChannelBusy_258(  )
       //.io_cyclesChannelBusy_257(  )
       //.io_cyclesChannelBusy_256(  )
       //.io_cyclesChannelBusy_255(  )
       //.io_cyclesChannelBusy_254(  )
       //.io_cyclesChannelBusy_253(  )
       //.io_cyclesChannelBusy_252(  )
       //.io_cyclesChannelBusy_251(  )
       //.io_cyclesChannelBusy_250(  )
       //.io_cyclesChannelBusy_249(  )
       //.io_cyclesChannelBusy_248(  )
       //.io_cyclesChannelBusy_247(  )
       //.io_cyclesChannelBusy_246(  )
       //.io_cyclesChannelBusy_245(  )
       //.io_cyclesChannelBusy_244(  )
       //.io_cyclesChannelBusy_243(  )
       //.io_cyclesChannelBusy_242(  )
       //.io_cyclesChannelBusy_241(  )
       //.io_cyclesChannelBusy_240(  )
       //.io_cyclesChannelBusy_239(  )
       //.io_cyclesChannelBusy_238(  )
       //.io_cyclesChannelBusy_237(  )
       //.io_cyclesChannelBusy_236(  )
       //.io_cyclesChannelBusy_235(  )
       //.io_cyclesChannelBusy_234(  )
       //.io_cyclesChannelBusy_233(  )
       //.io_cyclesChannelBusy_232(  )
       //.io_cyclesChannelBusy_231(  )
       //.io_cyclesChannelBusy_230(  )
       //.io_cyclesChannelBusy_229(  )
       //.io_cyclesChannelBusy_228(  )
       //.io_cyclesChannelBusy_227(  )
       //.io_cyclesChannelBusy_226(  )
       //.io_cyclesChannelBusy_225(  )
       //.io_cyclesChannelBusy_224(  )
       //.io_cyclesChannelBusy_223(  )
       //.io_cyclesChannelBusy_222(  )
       //.io_cyclesChannelBusy_221(  )
       //.io_cyclesChannelBusy_220(  )
       //.io_cyclesChannelBusy_219(  )
       //.io_cyclesChannelBusy_218(  )
       //.io_cyclesChannelBusy_217(  )
       //.io_cyclesChannelBusy_216(  )
       //.io_cyclesChannelBusy_215(  )
       //.io_cyclesChannelBusy_214(  )
       //.io_cyclesChannelBusy_213(  )
       //.io_cyclesChannelBusy_212(  )
       //.io_cyclesChannelBusy_211(  )
       //.io_cyclesChannelBusy_210(  )
       //.io_cyclesChannelBusy_209(  )
       //.io_cyclesChannelBusy_208(  )
       //.io_cyclesChannelBusy_207(  )
       //.io_cyclesChannelBusy_206(  )
       //.io_cyclesChannelBusy_205(  )
       //.io_cyclesChannelBusy_204(  )
       //.io_cyclesChannelBusy_203(  )
       //.io_cyclesChannelBusy_202(  )
       //.io_cyclesChannelBusy_201(  )
       //.io_cyclesChannelBusy_200(  )
       //.io_cyclesChannelBusy_199(  )
       //.io_cyclesChannelBusy_198(  )
       //.io_cyclesChannelBusy_197(  )
       //.io_cyclesChannelBusy_196(  )
       //.io_cyclesChannelBusy_195(  )
       //.io_cyclesChannelBusy_194(  )
       //.io_cyclesChannelBusy_193(  )
       //.io_cyclesChannelBusy_192(  )
       //.io_cyclesChannelBusy_191(  )
       //.io_cyclesChannelBusy_190(  )
       //.io_cyclesChannelBusy_189(  )
       //.io_cyclesChannelBusy_188(  )
       //.io_cyclesChannelBusy_187(  )
       //.io_cyclesChannelBusy_186(  )
       //.io_cyclesChannelBusy_185(  )
       //.io_cyclesChannelBusy_184(  )
       //.io_cyclesChannelBusy_183(  )
       //.io_cyclesChannelBusy_182(  )
       //.io_cyclesChannelBusy_181(  )
       //.io_cyclesChannelBusy_180(  )
       //.io_cyclesChannelBusy_179(  )
       //.io_cyclesChannelBusy_178(  )
       //.io_cyclesChannelBusy_177(  )
       //.io_cyclesChannelBusy_176(  )
       //.io_cyclesChannelBusy_175(  )
       //.io_cyclesChannelBusy_174(  )
       //.io_cyclesChannelBusy_173(  )
       //.io_cyclesChannelBusy_172(  )
       //.io_cyclesChannelBusy_171(  )
       //.io_cyclesChannelBusy_170(  )
       //.io_cyclesChannelBusy_169(  )
       //.io_cyclesChannelBusy_168(  )
       //.io_cyclesChannelBusy_167(  )
       //.io_cyclesChannelBusy_166(  )
       //.io_cyclesChannelBusy_165(  )
       //.io_cyclesChannelBusy_164(  )
       //.io_cyclesChannelBusy_163(  )
       //.io_cyclesChannelBusy_162(  )
       //.io_cyclesChannelBusy_161(  )
       //.io_cyclesChannelBusy_160(  )
       //.io_cyclesChannelBusy_159(  )
       //.io_cyclesChannelBusy_158(  )
       //.io_cyclesChannelBusy_157(  )
       //.io_cyclesChannelBusy_156(  )
       //.io_cyclesChannelBusy_155(  )
       //.io_cyclesChannelBusy_154(  )
       //.io_cyclesChannelBusy_153(  )
       //.io_cyclesChannelBusy_152(  )
       //.io_cyclesChannelBusy_151(  )
       //.io_cyclesChannelBusy_150(  )
       //.io_cyclesChannelBusy_149(  )
       //.io_cyclesChannelBusy_148(  )
       //.io_cyclesChannelBusy_147(  )
       //.io_cyclesChannelBusy_146(  )
       //.io_cyclesChannelBusy_145(  )
       //.io_cyclesChannelBusy_144(  )
       //.io_cyclesChannelBusy_143(  )
       //.io_cyclesChannelBusy_142(  )
       //.io_cyclesChannelBusy_141(  )
       //.io_cyclesChannelBusy_140(  )
       //.io_cyclesChannelBusy_139(  )
       //.io_cyclesChannelBusy_138(  )
       //.io_cyclesChannelBusy_137(  )
       //.io_cyclesChannelBusy_136(  )
       //.io_cyclesChannelBusy_135(  )
       //.io_cyclesChannelBusy_134(  )
       //.io_cyclesChannelBusy_133(  )
       //.io_cyclesChannelBusy_132(  )
       //.io_cyclesChannelBusy_131(  )
       //.io_cyclesChannelBusy_130(  )
       //.io_cyclesChannelBusy_129(  )
       //.io_cyclesChannelBusy_128(  )
       //.io_cyclesChannelBusy_127(  )
       //.io_cyclesChannelBusy_126(  )
       //.io_cyclesChannelBusy_125(  )
       //.io_cyclesChannelBusy_124(  )
       //.io_cyclesChannelBusy_123(  )
       //.io_cyclesChannelBusy_122(  )
       //.io_cyclesChannelBusy_121(  )
       //.io_cyclesChannelBusy_120(  )
       //.io_cyclesChannelBusy_119(  )
       //.io_cyclesChannelBusy_118(  )
       //.io_cyclesChannelBusy_117(  )
       //.io_cyclesChannelBusy_116(  )
       //.io_cyclesChannelBusy_115(  )
       //.io_cyclesChannelBusy_114(  )
       //.io_cyclesChannelBusy_113(  )
       //.io_cyclesChannelBusy_112(  )
       //.io_cyclesChannelBusy_111(  )
       //.io_cyclesChannelBusy_110(  )
       //.io_cyclesChannelBusy_109(  )
       //.io_cyclesChannelBusy_108(  )
       //.io_cyclesChannelBusy_107(  )
       //.io_cyclesChannelBusy_106(  )
       //.io_cyclesChannelBusy_105(  )
       //.io_cyclesChannelBusy_104(  )
       //.io_cyclesChannelBusy_103(  )
       //.io_cyclesChannelBusy_102(  )
       //.io_cyclesChannelBusy_101(  )
       //.io_cyclesChannelBusy_100(  )
       //.io_cyclesChannelBusy_99(  )
       //.io_cyclesChannelBusy_98(  )
       //.io_cyclesChannelBusy_97(  )
       //.io_cyclesChannelBusy_96(  )
       //.io_cyclesChannelBusy_95(  )
       //.io_cyclesChannelBusy_94(  )
       //.io_cyclesChannelBusy_93(  )
       //.io_cyclesChannelBusy_92(  )
       //.io_cyclesChannelBusy_91(  )
       //.io_cyclesChannelBusy_90(  )
       //.io_cyclesChannelBusy_89(  )
       //.io_cyclesChannelBusy_88(  )
       //.io_cyclesChannelBusy_87(  )
       //.io_cyclesChannelBusy_86(  )
       //.io_cyclesChannelBusy_85(  )
       //.io_cyclesChannelBusy_84(  )
       //.io_cyclesChannelBusy_83(  )
       //.io_cyclesChannelBusy_82(  )
       //.io_cyclesChannelBusy_81(  )
       //.io_cyclesChannelBusy_80(  )
       //.io_cyclesChannelBusy_79(  )
       //.io_cyclesChannelBusy_78(  )
       //.io_cyclesChannelBusy_77(  )
       //.io_cyclesChannelBusy_76(  )
       //.io_cyclesChannelBusy_75(  )
       //.io_cyclesChannelBusy_74(  )
       //.io_cyclesChannelBusy_73(  )
       //.io_cyclesChannelBusy_72(  )
       //.io_cyclesChannelBusy_71(  )
       //.io_cyclesChannelBusy_70(  )
       //.io_cyclesChannelBusy_69(  )
       //.io_cyclesChannelBusy_68(  )
       //.io_cyclesChannelBusy_67(  )
       //.io_cyclesChannelBusy_66(  )
       //.io_cyclesChannelBusy_65(  )
       //.io_cyclesChannelBusy_64(  )
       //.io_cyclesChannelBusy_63(  )
       //.io_cyclesChannelBusy_62(  )
       //.io_cyclesChannelBusy_61(  )
       //.io_cyclesChannelBusy_60(  )
       //.io_cyclesChannelBusy_59(  )
       //.io_cyclesChannelBusy_58(  )
       //.io_cyclesChannelBusy_57(  )
       //.io_cyclesChannelBusy_56(  )
       //.io_cyclesChannelBusy_55(  )
       //.io_cyclesChannelBusy_54(  )
       //.io_cyclesChannelBusy_53(  )
       //.io_cyclesChannelBusy_52(  )
       //.io_cyclesChannelBusy_51(  )
       //.io_cyclesChannelBusy_50(  )
       //.io_cyclesChannelBusy_49(  )
       //.io_cyclesChannelBusy_48(  )
       //.io_cyclesChannelBusy_47(  )
       //.io_cyclesChannelBusy_46(  )
       //.io_cyclesChannelBusy_45(  )
       //.io_cyclesChannelBusy_44(  )
       //.io_cyclesChannelBusy_43(  )
       //.io_cyclesChannelBusy_42(  )
       //.io_cyclesChannelBusy_41(  )
       //.io_cyclesChannelBusy_40(  )
       //.io_cyclesChannelBusy_39(  )
       //.io_cyclesChannelBusy_38(  )
       //.io_cyclesChannelBusy_37(  )
       //.io_cyclesChannelBusy_36(  )
       //.io_cyclesChannelBusy_35(  )
       //.io_cyclesChannelBusy_34(  )
       //.io_cyclesChannelBusy_33(  )
       //.io_cyclesChannelBusy_32(  )
       //.io_cyclesChannelBusy_31(  )
       //.io_cyclesChannelBusy_30(  )
       //.io_cyclesChannelBusy_29(  )
       //.io_cyclesChannelBusy_28(  )
       //.io_cyclesChannelBusy_27(  )
       //.io_cyclesChannelBusy_26(  )
       //.io_cyclesChannelBusy_25(  )
       //.io_cyclesChannelBusy_24(  )
       //.io_cyclesChannelBusy_23(  )
       //.io_cyclesChannelBusy_22(  )
       //.io_cyclesChannelBusy_21(  )
       //.io_cyclesChannelBusy_20(  )
       //.io_cyclesChannelBusy_19(  )
       //.io_cyclesChannelBusy_18(  )
       //.io_cyclesChannelBusy_17(  )
       //.io_cyclesChannelBusy_16(  )
       //.io_cyclesChannelBusy_15(  )
       .io_cyclesChannelBusy_14( VCCMesh_io_cyclesChannelBusy_14 ),
       .io_cyclesChannelBusy_13( VCCMesh_io_cyclesChannelBusy_13 ),
       .io_cyclesChannelBusy_12( VCCMesh_io_cyclesChannelBusy_12 ),
       .io_cyclesChannelBusy_11( VCCMesh_io_cyclesChannelBusy_11 ),
       .io_cyclesChannelBusy_10( VCCMesh_io_cyclesChannelBusy_10 ),
       .io_cyclesChannelBusy_9( VCCMesh_io_cyclesChannelBusy_9 ),
       .io_cyclesChannelBusy_8( VCCMesh_io_cyclesChannelBusy_8 ),
       .io_cyclesChannelBusy_7( VCCMesh_io_cyclesChannelBusy_7 ),
       .io_cyclesChannelBusy_6( VCCMesh_io_cyclesChannelBusy_6 ),
       .io_cyclesChannelBusy_5( VCCMesh_io_cyclesChannelBusy_5 ),
       .io_cyclesChannelBusy_4( VCCMesh_io_cyclesChannelBusy_4 ),
       .io_cyclesChannelBusy_3( VCCMesh_io_cyclesChannelBusy_3 ),
       .io_cyclesChannelBusy_2( VCCMesh_io_cyclesChannelBusy_2 ),
       .io_cyclesChannelBusy_1( VCCMesh_io_cyclesChannelBusy_1 ),
       .io_cyclesChannelBusy_0( VCCMesh_io_cyclesChannelBusy_0 ),
       .io_bypass_2( io_bypass_2 ),
       .io_bypass_1( io_bypass_1 ),
       .io_bypass_0( io_bypass_0 )
  );
`ifndef SYNTHESIS
// synthesis translate_off
    assign VCCMesh.io_cyclesChannelBusy_14 = {1{1'b0}};
    assign VCCMesh.io_cyclesChannelBusy_13 = {1{1'b0}};
    assign VCCMesh.io_cyclesChannelBusy_11 = {1{1'b0}};
    assign VCCMesh.io_cyclesChannelBusy_10 = {1{1'b0}};
    assign VCCMesh.io_cyclesChannelBusy_9 = {1{1'b0}};
    assign VCCMesh.io_cyclesChannelBusy_8 = {1{1'b0}};
    assign VCCMesh.io_cyclesChannelBusy_5 = {1{1'b0}};
    assign VCCMesh.io_cyclesChannelBusy_4 = {1{1'b0}};
    assign VCCMesh.io_cyclesChannelBusy_3 = {1{1'b0}};
    assign VCCMesh.io_cyclesChannelBusy_2 = {1{1'b0}};
    assign VCCMesh.io_cyclesChannelBusy_0 = {1{1'b0}};
// synthesis translate_on
`endif
  InjectionChannelQ InjectionChannelQ(.clk(clk), .reset(reset),
       .io_in_flit_x( InputPacketInterface_io_out_flit_x ),
       .io_in_flitValid( InputPacketInterface_io_out_flitValid ),
       .io_in_credit_grant( InjectionChannelQ_io_in_credit_grant ),
       .io_out_flit_x( InjectionChannelQ_io_out_flit_x ),
       .io_out_flitValid( InjectionChannelQ_io_out_flitValid ),
       .io_out_credit_1_grant( VCCMesh_io_inChannels_0_credit_1_grant ),
       .io_out_credit_0_grant( VCCMesh_io_inChannels_0_credit_0_grant )
  );
  EjectionChannelQ EjectionChannelQ(.clk(clk), .reset(reset),
       .io_in_flit_x( VCCMesh_io_outChannels_0_flit_x ),
       .io_in_flitValid( VCCMesh_io_outChannels_0_flitValid ),
       .io_in_credit_1_grant( EjectionChannelQ_io_in_credit_1_grant ),
       .io_in_credit_0_grant( EjectionChannelQ_io_in_credit_0_grant ),
       .io_out_flit_x( EjectionChannelQ_io_out_flit_x ),
       .io_out_flitValid( EjectionChannelQ_io_out_flitValid ),
       .io_out_credit_grant( io_ports_0_out_credit_grant )
  );
  InputPacketInterface InputPacketInterface(.clk(clk), .reset(reset),
       .io_in_ready( InputPacketInterface_io_in_ready ),
       .io_in_valid( io_ports_0_in_packetValid ),
       .io_in_bits_x( io_ports_0_in_packet_x ),
       .io_out_flit_x( InputPacketInterface_io_out_flit_x ),
       .io_out_flitValid( InputPacketInterface_io_out_flitValid ),
       .io_out_credit_grant( InjectionChannelQ_io_in_credit_grant )
  );
  InjectionChannelQ InjectionChannelQ_1(.clk(clk), .reset(reset),
       .io_in_flit_x( InputPacketInterface_1_io_out_flit_x ),
       .io_in_flitValid( InputPacketInterface_1_io_out_flitValid ),
       .io_in_credit_grant( InjectionChannelQ_1_io_in_credit_grant ),
       .io_out_flit_x( InjectionChannelQ_1_io_out_flit_x ),
       .io_out_flitValid( InjectionChannelQ_1_io_out_flitValid ),
       .io_out_credit_1_grant( VCCMesh_io_inChannels_1_credit_1_grant ),
       .io_out_credit_0_grant( VCCMesh_io_inChannels_1_credit_0_grant )
  );
  EjectionChannelQ EjectionChannelQ_1(.clk(clk), .reset(reset),
       .io_in_flit_x( VCCMesh_io_outChannels_1_flit_x ),
       .io_in_flitValid( VCCMesh_io_outChannels_1_flitValid ),
       .io_in_credit_1_grant( EjectionChannelQ_1_io_in_credit_1_grant ),
       .io_in_credit_0_grant( EjectionChannelQ_1_io_in_credit_0_grant ),
       .io_out_flit_x( EjectionChannelQ_1_io_out_flit_x ),
       .io_out_flitValid( EjectionChannelQ_1_io_out_flitValid ),
       .io_out_credit_grant( io_ports_1_out_credit_grant )
  );
  InputPacketInterface InputPacketInterface_1(.clk(clk), .reset(reset),
       .io_in_ready( InputPacketInterface_1_io_in_ready ),
       .io_in_valid( io_ports_1_in_packetValid ),
       .io_in_bits_x( io_ports_1_in_packet_x ),
       .io_out_flit_x( InputPacketInterface_1_io_out_flit_x ),
       .io_out_flitValid( InputPacketInterface_1_io_out_flitValid ),
       .io_out_credit_grant( InjectionChannelQ_1_io_in_credit_grant )
  );
  InjectionChannelQ InjectionChannelQ_2(.clk(clk), .reset(reset),
       .io_in_flit_x( InputPacketInterface_2_io_out_flit_x ),
       .io_in_flitValid( InputPacketInterface_2_io_out_flitValid ),
       .io_in_credit_grant( InjectionChannelQ_2_io_in_credit_grant ),
       .io_out_flit_x( InjectionChannelQ_2_io_out_flit_x ),
       .io_out_flitValid( InjectionChannelQ_2_io_out_flitValid ),
       .io_out_credit_1_grant( VCCMesh_io_inChannels_2_credit_1_grant ),
       .io_out_credit_0_grant( VCCMesh_io_inChannels_2_credit_0_grant )
  );
  EjectionChannelQ EjectionChannelQ_2(.clk(clk), .reset(reset),
       .io_in_flit_x( VCCMesh_io_outChannels_2_flit_x ),
       .io_in_flitValid( VCCMesh_io_outChannels_2_flitValid ),
       .io_in_credit_1_grant( EjectionChannelQ_2_io_in_credit_1_grant ),
       .io_in_credit_0_grant( EjectionChannelQ_2_io_in_credit_0_grant ),
       .io_out_flit_x( EjectionChannelQ_2_io_out_flit_x ),
       .io_out_flitValid( EjectionChannelQ_2_io_out_flitValid ),
       .io_out_credit_grant( io_ports_2_out_credit_grant )
  );
  InputPacketInterface InputPacketInterface_2(.clk(clk), .reset(reset),
       .io_in_ready( InputPacketInterface_2_io_in_ready ),
       .io_in_valid( io_ports_2_in_packetValid ),
       .io_in_bits_x( io_ports_2_in_packet_x ),
       .io_out_flit_x( InputPacketInterface_2_io_out_flit_x ),
       .io_out_flitValid( InputPacketInterface_2_io_out_flitValid ),
       .io_out_credit_grant( InjectionChannelQ_2_io_in_credit_grant )
  );
endmodule

module HeadBundle2Flit(
    input [15:0] io_inHead_packetID,
    input  io_inHead_isTail,
    input  io_inHead_vcPort,
    input [3:0] io_inHead_packetType,
    input [1:0] io_inHead_destination_2,
    input [1:0] io_inHead_destination_1,
    input [1:0] io_inHead_destination_0,
    input [2:0] io_inHead_priorityLevel,
    output[54:0] io_outFlit_x
);

  wire[54:0] T0;
  wire[54:0] T1;
  wire[31:0] T2;
  wire[30:0] T3;
  wire[30:0] T4;
  wire[8:0] T5;
  wire[4:0] T6;
  wire[3:0] T7;
  wire[21:0] T8;
  wire[4:0] T9;
  wire[16:0] T10;


  assign io_outFlit_x = T0;
  assign T0 = T1;
  assign T1 = {23'h0, T2};
  assign T2 = {T3, 1'h1};
  assign T3 = T4;
  assign T4 = {T8, T5};
  assign T5 = {T7, T6};
  assign T6 = {io_inHead_destination_0, io_inHead_priorityLevel};
  assign T7 = {io_inHead_destination_2, io_inHead_destination_1};
  assign T8 = {T10, T9};
  assign T9 = {io_inHead_vcPort, io_inHead_packetType};
  assign T10 = {io_inHead_packetID, io_inHead_isTail};
endmodule

module BodyBundle2Flit(
    input [15:0] io_inBody_packetID,
    input  io_inBody_isTail,
    input  io_inBody_vcPort,
    input [3:0] io_inBody_flitID,
    input [31:0] io_inBody_payload,
    output[54:0] io_outFlit_x
);

  wire[54:0] T0;
  wire[54:0] T1;
  wire[53:0] T2;
  wire[53:0] T3;
  wire[36:0] T4;
  wire[35:0] T5;
  wire[16:0] T6;


  assign io_outFlit_x = T0;
  assign T0 = T1;
  assign T1 = {T2, 1'h0};
  assign T2 = T3;
  assign T3 = {T6, T4};
  assign T4 = {io_inBody_vcPort, T5};
  assign T5 = {io_inBody_flitID, io_inBody_payload};
  assign T6 = {io_inBody_packetID, io_inBody_isTail};
endmodule

module PortDataGen(input clk, input reset,
    output io_config_ready,
    input  io_config_valid,
    input  io_config_bits_sequence,
    input [1:0] io_config_bits_destination_2,
    input [1:0] io_config_bits_destination_1,
    input [1:0] io_config_bits_destination_0,
    input [31:0] io_config_bits_count,
    output[54:0] io_out_packet_x,
    input  io_out_packetReady,
    output io_out_packetValid
);

  wire[31:0] T0;
  wire[31:0] T1;
  reg [15:0] lfsr;
  wire[15:0] T70;
  wire[15:0] T2;
  wire[14:0] T3;
  wire T4;
  wire T5;
  wire T6;
  wire T7;
  wire T8;
  wire T9;
  wire T10;
  wire[15:0] T11;
  reg [15:0] lfsr_prev;
  wire[15:0] T71;
  reg [31:0] count;
  wire[31:0] T72;
  wire[31:0] T12;
  wire[31:0] T13;
  wire T14;
  wire T15;
  wire T16;
  reg [1:0] state;
  wire[1:0] T73;
  wire[1:0] T17;
  wire[1:0] T18;
  wire[1:0] T19;
  wire[1:0] T20;
  wire[1:0] T21;
  wire T22;
  wire T23;
  wire T24;
  reg [6:0] initCount;
  wire[6:0] T74;
  wire[6:0] T25;
  wire[6:0] T26;
  wire T27;
  wire T28;
  wire T29;
  wire T30;
  wire T31;
  reg [31:0] config_count;
  wire[31:0] T32;
  wire[31:0] T33;
  wire T34;
  wire T35;
  wire[31:0] T36;
  wire T37;
  wire T38;
  wire T39;
  wire T40;
  wire T41;
  wire T42;
  wire T43;
  wire T44;
  wire T45;
  wire T46;
  wire[31:0] T47;
  wire T48;
  wire T49;
  wire T50;
  wire T51;
  reg  config_sequence;
  wire T52;
  reg  flip;
  wire T53;
  wire T54;
  reg [1:0] config_destination_0;
  wire[1:0] T55;
  reg [1:0] config_destination_1;
  wire[1:0] T56;
  reg [1:0] config_destination_2;
  wire[1:0] T57;
  wire T58;
  wire T59;
  wire T60;
  wire T61;
  wire[54:0] T62;
  wire[54:0] T63;
  wire[54:0] T64;
  wire[54:0] T65;
  wire T66;
  wire T67;
  wire T68;
  wire T69;
  wire[54:0] headExtract_io_outFlit_x;
  wire[54:0] bodyExtract_io_outFlit_x;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    lfsr = {1{1'b0}};
    lfsr_prev = {1{1'b0}};
    count = {1{1'b0}};
    state = {1{1'b0}};
    initCount = {1{1'b0}};
    config_count = {1{1'b0}};
    config_sequence = {1{1'b0}};
    flip = {1{1'b0}};
    config_destination_0 = {1{1'b0}};
    config_destination_1 = {1{1'b0}};
    config_destination_2 = {1{1'b0}};
  end
// synthesis translate_on
`endif

  assign T0 = config_sequence ? count : T1;
  assign T1 = {T11, lfsr};
  assign T70 = reset ? 16'h1 : T2;
  assign T2 = {T4, T3};
  assign T3 = lfsr[4'hf:1'h1];
  assign T4 = T6 ^ T5;
  assign T5 = lfsr[3'h5:3'h5];
  assign T6 = T8 ^ T7;
  assign T7 = lfsr[2'h3:2'h3];
  assign T8 = T10 ^ T9;
  assign T9 = lfsr[2'h2:2'h2];
  assign T10 = lfsr[1'h0:1'h0];
  assign T11 = lfsr ^ lfsr_prev;
  assign T71 = reset ? 16'hf25a : lfsr;
  assign T72 = reset ? 32'ha : T12;
  assign T12 = T14 ? T13 : count;
  assign T13 = count + 32'h1;
  assign T14 = T15 & io_out_packetReady;
  assign T15 = T50 & T16;
  assign T16 = state == 2'h3;
  assign T73 = reset ? 2'h0 : T17;
  assign T17 = T48 ? 2'h2 : T18;
  assign T18 = T45 ? 2'h1 : T19;
  assign T19 = T40 ? 2'h3 : T20;
  assign T20 = T29 ? 2'h2 : T21;
  assign T21 = T22 ? 2'h1 : state;
  assign T22 = T28 & T23;
  assign T23 = T24 ^ 1'h1;
  assign T24 = initCount != 7'h0;
  assign T74 = reset ? 7'h40 : T25;
  assign T25 = T27 ? T26 : initCount;
  assign T26 = initCount - 7'h1;
  assign T27 = T28 & T24;
  assign T28 = state == 2'h0;
  assign T29 = T37 & T30;
  assign T30 = T31 ^ 1'h1;
  assign T31 = config_count == 32'h0;
  assign T32 = T14 ? T36 : T33;
  assign T33 = T34 ? io_config_bits_count : config_count;
  assign T34 = T35 & io_config_valid;
  assign T35 = T37 & T31;
  assign T36 = config_count - 32'h1;
  assign T37 = T39 & T38;
  assign T38 = state == 2'h1;
  assign T39 = T28 ^ 1'h1;
  assign T40 = T41 & io_out_packetReady;
  assign T41 = T43 & T42;
  assign T42 = state == 2'h2;
  assign T43 = T44 ^ 1'h1;
  assign T44 = T28 | T38;
  assign T45 = T14 & T46;
  assign T46 = T47 == 32'h0;
  assign T47 = config_count - 32'h1;
  assign T48 = T14 & T49;
  assign T49 = T46 ^ 1'h1;
  assign T50 = T51 ^ 1'h1;
  assign T51 = T44 | T42;
  assign T52 = T34 ? io_config_bits_sequence : config_sequence;
  assign T53 = T14 ? T54 : flip;
  assign T54 = ~ flip;
  assign T55 = T34 ? io_config_bits_destination_0 : config_destination_0;
  assign T56 = T34 ? io_config_bits_destination_1 : config_destination_1;
  assign T57 = T34 ? io_config_bits_destination_2 : config_destination_2;
  assign io_out_packetValid = T58;
  assign T58 = T14 ? 1'h1 : T59;
  assign T59 = T40 ? 1'h1 : T60;
  assign T60 = T37 ? 1'h0 : T61;
  assign T61 = T28 ? 1'h0 : 1'h0;
  assign io_out_packet_x = T62;
  assign T62 = T14 ? bodyExtract_io_outFlit_x : T63;
  assign T63 = T40 ? headExtract_io_outFlit_x : T64;
  assign T64 = T37 ? 55'h0 : T65;
  assign T65 = T28 ? 55'h0 : 55'h0;
  assign io_config_ready = T66;
  assign T66 = T15 ? 1'h0 : T67;
  assign T67 = T41 ? 1'h0 : T68;
  assign T68 = T35 ? 1'h1 : T69;
  assign T69 = T28 ? 1'h0 : 1'h0;
  HeadBundle2Flit headExtract(
       .io_inHead_packetID( 16'h0 ),
       .io_inHead_isTail( 1'h0 ),
       .io_inHead_vcPort( flip ),
       .io_inHead_packetType( 4'h0 ),
       .io_inHead_destination_2( config_destination_2 ),
       .io_inHead_destination_1( config_destination_1 ),
       .io_inHead_destination_0( config_destination_0 ),
       .io_inHead_priorityLevel( 3'h0 ),
       .io_outFlit_x( headExtract_io_outFlit_x )
  );
  BodyBundle2Flit bodyExtract(
       .io_inBody_packetID( 16'h0 ),
       .io_inBody_isTail( 1'h1 ),
       .io_inBody_vcPort( flip ),
       .io_inBody_flitID( 4'h0 ),
       .io_inBody_payload( T0 ),
       .io_outFlit_x( bodyExtract_io_outFlit_x )
  );

  always @(posedge clk) begin
    if(reset) begin
      lfsr <= 16'h1;
    end else begin
      lfsr <= T2;
    end
    if(reset) begin
      lfsr_prev <= 16'hf25a;
    end else begin
      lfsr_prev <= lfsr;
    end
    if(reset) begin
      count <= 32'ha;
    end else if(T14) begin
      count <= T13;
    end
    if(reset) begin
      state <= 2'h0;
    end else if(T48) begin
      state <= 2'h2;
    end else if(T45) begin
      state <= 2'h1;
    end else if(T40) begin
      state <= 2'h3;
    end else if(T29) begin
      state <= 2'h2;
    end else if(T22) begin
      state <= 2'h1;
    end
    if(reset) begin
      initCount <= 7'h40;
    end else if(T27) begin
      initCount <= T26;
    end
    if(T14) begin
      config_count <= T36;
    end else if(T34) begin
      config_count <= io_config_bits_count;
    end
    if(T34) begin
      config_sequence <= io_config_bits_sequence;
    end
    if(T14) begin
      flip <= T54;
    end
    if(T34) begin
      config_destination_0 <= io_config_bits_destination_0;
    end
    if(T34) begin
      config_destination_1 <= io_config_bits_destination_1;
    end
    if(T34) begin
      config_destination_2 <= io_config_bits_destination_2;
    end
  end
endmodule

module PortDataSink(input clk, input reset,
    input [54:0] io_in_flit_x,
    input  io_in_flitValid,
    output io_in_credit_grant,
    output[31:0] io_count,
    output[54:0] io_dump
);

  reg [54:0] dump;
  wire[54:0] T0;
  wire[54:0] T1;
  wire[54:0] T2;
  reg [31:0] count;
  wire[31:0] T5;
  wire[31:0] T3;
  wire[31:0] T4;

`ifndef SYNTHESIS
// synthesis translate_off
  integer initvar;
  initial begin
    #0.002;
    dump = {2{1'b0}};
    count = {1{1'b0}};
  end
// synthesis translate_on
`endif

  assign io_dump = dump;
  assign T0 = io_in_flitValid ? T1 : dump;
  assign T1 = dump ^ T2;
  assign T2 = io_in_flit_x;
  assign io_count = count;
  assign T5 = reset ? 32'h0 : T3;
  assign T3 = io_in_flitValid ? T4 : count;
  assign T4 = count + 32'h1;
  assign io_in_credit_grant = 1'h1;

  always @(posedge clk) begin
    if(io_in_flitValid) begin
      dump <= T1;
    end
    if(reset) begin
      count <= 32'h0;
    end else if(io_in_flitValid) begin
      count <= T4;
    end
  end
endmodule

module My_MeshWrapper(input clk, input reset,
    output io_config_2_ready,
    input  io_config_2_valid,
    input  io_config_2_bits_sequence,
    input [1:0] io_config_2_bits_destination_2,
    input [1:0] io_config_2_bits_destination_1,
    input [1:0] io_config_2_bits_destination_0,
    input [31:0] io_config_2_bits_count,
    output io_config_1_ready,
    input  io_config_1_valid,
    input  io_config_1_bits_sequence,
    input [1:0] io_config_1_bits_destination_2,
    input [1:0] io_config_1_bits_destination_1,
    input [1:0] io_config_1_bits_destination_0,
    input [31:0] io_config_1_bits_count,
    output io_config_0_ready,
    input  io_config_0_valid,
    input  io_config_0_bits_sequence,
    input [1:0] io_config_0_bits_destination_2,
    input [1:0] io_config_0_bits_destination_1,
    input [1:0] io_config_0_bits_destination_0,
    input [31:0] io_config_0_bits_count,
    output[31:0] io_count_2,
    output[31:0] io_count_1,
    output[31:0] io_count_0,
    output[54:0] io_dump_2,
    output[54:0] io_dump_1,
    output[54:0] io_dump_0,
    input  io_bypass_2,
    input  io_bypass_1,
    input  io_bypass_0
);

  wire PortDataSink_io_in_credit_grant;
  wire[31:0] PortDataSink_io_count;
  wire[54:0] PortDataSink_io_dump;
  wire PortDataSink_1_io_in_credit_grant;
  wire[31:0] PortDataSink_1_io_count;
  wire[54:0] PortDataSink_1_io_dump;
  wire PortDataSink_2_io_in_credit_grant;
  wire[31:0] PortDataSink_2_io_count;
  wire[54:0] PortDataSink_2_io_dump;
  wire PortDataGen_io_config_ready;
  wire[54:0] PortDataGen_io_out_packet_x;
  wire PortDataGen_io_out_packetValid;
  wire PortDataGen_1_io_config_ready;
  wire[54:0] PortDataGen_1_io_out_packet_x;
  wire PortDataGen_1_io_out_packetValid;
  wire PortDataGen_2_io_config_ready;
  wire[54:0] PortDataGen_2_io_out_packet_x;
  wire PortDataGen_2_io_out_packetValid;
  wire mesh_io_ports_2_in_packetReady;
  wire[54:0] mesh_io_ports_2_out_flit_x;
  wire mesh_io_ports_2_out_flitValid;
  wire mesh_io_ports_1_in_packetReady;
  wire[54:0] mesh_io_ports_1_out_flit_x;
  wire mesh_io_ports_1_out_flitValid;
  wire mesh_io_ports_0_in_packetReady;
  wire[54:0] mesh_io_ports_0_out_flit_x;
  wire mesh_io_ports_0_out_flitValid;


  assign io_dump_0 = PortDataSink_io_dump;
  assign io_dump_1 = PortDataSink_1_io_dump;
  assign io_dump_2 = PortDataSink_2_io_dump;
  assign io_count_0 = PortDataSink_io_count;
  assign io_count_1 = PortDataSink_1_io_count;
  assign io_count_2 = PortDataSink_2_io_count;
  assign io_config_0_ready = PortDataGen_io_config_ready;
  assign io_config_1_ready = PortDataGen_1_io_config_ready;
  assign io_config_2_ready = PortDataGen_2_io_config_ready;
  My_Mesh mesh(.clk(clk), .reset(reset),
       .io_ports_2_in_packet_x( PortDataGen_2_io_out_packet_x ),
       .io_ports_2_in_packetReady( mesh_io_ports_2_in_packetReady ),
       .io_ports_2_in_packetValid( PortDataGen_2_io_out_packetValid ),
       .io_ports_2_out_flit_x( mesh_io_ports_2_out_flit_x ),
       .io_ports_2_out_flitValid( mesh_io_ports_2_out_flitValid ),
       .io_ports_2_out_credit_grant( PortDataSink_2_io_in_credit_grant ),
       .io_ports_1_in_packet_x( PortDataGen_1_io_out_packet_x ),
       .io_ports_1_in_packetReady( mesh_io_ports_1_in_packetReady ),
       .io_ports_1_in_packetValid( PortDataGen_1_io_out_packetValid ),
       .io_ports_1_out_flit_x( mesh_io_ports_1_out_flit_x ),
       .io_ports_1_out_flitValid( mesh_io_ports_1_out_flitValid ),
       .io_ports_1_out_credit_grant( PortDataSink_1_io_in_credit_grant ),
       .io_ports_0_in_packet_x( PortDataGen_io_out_packet_x ),
       .io_ports_0_in_packetReady( mesh_io_ports_0_in_packetReady ),
       .io_ports_0_in_packetValid( PortDataGen_io_out_packetValid ),
       .io_ports_0_out_flit_x( mesh_io_ports_0_out_flit_x ),
       .io_ports_0_out_flitValid( mesh_io_ports_0_out_flitValid ),
       .io_ports_0_out_credit_grant( PortDataSink_io_in_credit_grant ),
       .io_bypass_2( io_bypass_2 ),
       .io_bypass_1( io_bypass_1 ),
       .io_bypass_0( io_bypass_0 )
       //.io_cyclesRouterBusy_2(  )
       //.io_cyclesRouterBusy_1(  )
       //.io_cyclesRouterBusy_0(  )
       //.io_cyclesChannelBusy_14(  )
       //.io_cyclesChannelBusy_13(  )
       //.io_cyclesChannelBusy_12(  )
       //.io_cyclesChannelBusy_11(  )
       //.io_cyclesChannelBusy_10(  )
       //.io_cyclesChannelBusy_9(  )
       //.io_cyclesChannelBusy_8(  )
       //.io_cyclesChannelBusy_7(  )
       //.io_cyclesChannelBusy_6(  )
       //.io_cyclesChannelBusy_5(  )
       //.io_cyclesChannelBusy_4(  )
       //.io_cyclesChannelBusy_3(  )
       //.io_cyclesChannelBusy_2(  )
       //.io_cyclesChannelBusy_1(  )
       //.io_cyclesChannelBusy_0(  )
  );
  PortDataGen PortDataGen(.clk(clk), .reset(reset),
       .io_config_ready( PortDataGen_io_config_ready ),
       .io_config_valid( io_config_0_valid ),
       .io_config_bits_sequence( io_config_0_bits_sequence ),
       .io_config_bits_destination_2( io_config_0_bits_destination_2 ),
       .io_config_bits_destination_1( io_config_0_bits_destination_1 ),
       .io_config_bits_destination_0( io_config_0_bits_destination_0 ),
       .io_config_bits_count( io_config_0_bits_count ),
       .io_out_packet_x( PortDataGen_io_out_packet_x ),
       .io_out_packetReady( mesh_io_ports_0_in_packetReady ),
       .io_out_packetValid( PortDataGen_io_out_packetValid )
  );
  PortDataGen PortDataGen_1(.clk(clk), .reset(reset),
       .io_config_ready( PortDataGen_1_io_config_ready ),
       .io_config_valid( io_config_1_valid ),
       .io_config_bits_sequence( io_config_1_bits_sequence ),
       .io_config_bits_destination_2( io_config_1_bits_destination_2 ),
       .io_config_bits_destination_1( io_config_1_bits_destination_1 ),
       .io_config_bits_destination_0( io_config_1_bits_destination_0 ),
       .io_config_bits_count( io_config_1_bits_count ),
       .io_out_packet_x( PortDataGen_1_io_out_packet_x ),
       .io_out_packetReady( mesh_io_ports_1_in_packetReady ),
       .io_out_packetValid( PortDataGen_1_io_out_packetValid )
  );
  PortDataGen PortDataGen_2(.clk(clk), .reset(reset),
       .io_config_ready( PortDataGen_2_io_config_ready ),
       .io_config_valid( io_config_2_valid ),
       .io_config_bits_sequence( io_config_2_bits_sequence ),
       .io_config_bits_destination_2( io_config_2_bits_destination_2 ),
       .io_config_bits_destination_1( io_config_2_bits_destination_1 ),
       .io_config_bits_destination_0( io_config_2_bits_destination_0 ),
       .io_config_bits_count( io_config_2_bits_count ),
       .io_out_packet_x( PortDataGen_2_io_out_packet_x ),
       .io_out_packetReady( mesh_io_ports_2_in_packetReady ),
       .io_out_packetValid( PortDataGen_2_io_out_packetValid )
  );
  PortDataSink PortDataSink(.clk(clk), .reset(reset),
       .io_in_flit_x( mesh_io_ports_0_out_flit_x ),
       .io_in_flitValid( mesh_io_ports_0_out_flitValid ),
       .io_in_credit_grant( PortDataSink_io_in_credit_grant ),
       .io_count( PortDataSink_io_count ),
       .io_dump( PortDataSink_io_dump )
  );
  PortDataSink PortDataSink_1(.clk(clk), .reset(reset),
       .io_in_flit_x( mesh_io_ports_1_out_flit_x ),
       .io_in_flitValid( mesh_io_ports_1_out_flitValid ),
       .io_in_credit_grant( PortDataSink_1_io_in_credit_grant ),
       .io_count( PortDataSink_1_io_count ),
       .io_dump( PortDataSink_1_io_dump )
  );
  PortDataSink PortDataSink_2(.clk(clk), .reset(reset),
       .io_in_flit_x( mesh_io_ports_2_out_flit_x ),
       .io_in_flitValid( mesh_io_ports_2_out_flitValid ),
       .io_in_credit_grant( PortDataSink_2_io_in_credit_grant ),
       .io_count( PortDataSink_2_io_count ),
       .io_dump( PortDataSink_2_io_dump )
  );
endmodule

